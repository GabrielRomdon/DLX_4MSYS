
module REG_GENERIC_NBIT32_0 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163;

  DFF_X1 \DATA_OUT_reg[17]  ( .D(n146), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n161), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n162), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n163), .CK(CLK), .Q(DATA_OUT[0]) );
  BUF_X1 U31 ( .A(n130), .Z(n93) );
  BUF_X1 U32 ( .A(n130), .Z(n94) );
  BUF_X1 U33 ( .A(n89), .Z(n90) );
  BUF_X1 U34 ( .A(n89), .Z(n91) );
  BUF_X2 U35 ( .A(n130), .Z(n95) );
  BUF_X1 U36 ( .A(n89), .Z(n92) );
  AND2_X1 U37 ( .A1(n96), .A2(n98), .ZN(n89) );
  INV_X1 U38 ( .A(n97), .ZN(n96) );
  INV_X1 U39 ( .A(RST), .ZN(n97) );
  OR2_X1 U40 ( .A1(EN), .A2(n97), .ZN(n98) );
  INV_X1 U41 ( .A(n98), .ZN(n130) );
  AOI22_X1 U42 ( .A1(DATA_OUT[0]), .A2(n93), .B1(DATA_IN[0]), .B2(n90), .ZN(
        n99) );
  INV_X1 U43 ( .A(n99), .ZN(n163) );
  AOI22_X1 U44 ( .A1(DATA_OUT[1]), .A2(n93), .B1(DATA_IN[1]), .B2(n90), .ZN(
        n100) );
  INV_X1 U45 ( .A(n100), .ZN(n162) );
  AOI22_X1 U46 ( .A1(DATA_OUT[2]), .A2(n93), .B1(DATA_IN[2]), .B2(n90), .ZN(
        n101) );
  INV_X1 U47 ( .A(n101), .ZN(n161) );
  AOI22_X1 U48 ( .A1(DATA_OUT[3]), .A2(n93), .B1(DATA_IN[3]), .B2(n90), .ZN(
        n102) );
  INV_X1 U49 ( .A(n102), .ZN(n160) );
  AOI22_X1 U50 ( .A1(DATA_OUT[4]), .A2(n93), .B1(DATA_IN[4]), .B2(n90), .ZN(
        n103) );
  INV_X1 U51 ( .A(n103), .ZN(n159) );
  AOI22_X1 U52 ( .A1(DATA_OUT[5]), .A2(n93), .B1(DATA_IN[5]), .B2(n90), .ZN(
        n104) );
  INV_X1 U53 ( .A(n104), .ZN(n158) );
  AOI22_X1 U54 ( .A1(DATA_OUT[6]), .A2(n93), .B1(DATA_IN[6]), .B2(n90), .ZN(
        n105) );
  INV_X1 U55 ( .A(n105), .ZN(n157) );
  AOI22_X1 U56 ( .A1(DATA_OUT[7]), .A2(n93), .B1(DATA_IN[7]), .B2(n90), .ZN(
        n106) );
  INV_X1 U57 ( .A(n106), .ZN(n156) );
  AOI22_X1 U58 ( .A1(DATA_OUT[8]), .A2(n93), .B1(DATA_IN[8]), .B2(n90), .ZN(
        n107) );
  INV_X1 U59 ( .A(n107), .ZN(n155) );
  AOI22_X1 U60 ( .A1(DATA_OUT[9]), .A2(n93), .B1(DATA_IN[9]), .B2(n90), .ZN(
        n108) );
  INV_X1 U61 ( .A(n108), .ZN(n154) );
  AOI22_X1 U62 ( .A1(DATA_OUT[10]), .A2(n93), .B1(DATA_IN[10]), .B2(n90), .ZN(
        n109) );
  INV_X1 U63 ( .A(n109), .ZN(n153) );
  AOI22_X1 U64 ( .A1(DATA_OUT[11]), .A2(n93), .B1(DATA_IN[11]), .B2(n90), .ZN(
        n110) );
  INV_X1 U65 ( .A(n110), .ZN(n152) );
  AOI22_X1 U66 ( .A1(DATA_OUT[12]), .A2(n94), .B1(DATA_IN[12]), .B2(n91), .ZN(
        n111) );
  INV_X1 U67 ( .A(n111), .ZN(n151) );
  AOI22_X1 U68 ( .A1(DATA_OUT[13]), .A2(n94), .B1(DATA_IN[13]), .B2(n91), .ZN(
        n112) );
  INV_X1 U69 ( .A(n112), .ZN(n150) );
  AOI22_X1 U70 ( .A1(DATA_OUT[14]), .A2(n94), .B1(DATA_IN[14]), .B2(n91), .ZN(
        n113) );
  INV_X1 U71 ( .A(n113), .ZN(n149) );
  AOI22_X1 U72 ( .A1(DATA_OUT[15]), .A2(n94), .B1(DATA_IN[15]), .B2(n91), .ZN(
        n114) );
  INV_X1 U73 ( .A(n114), .ZN(n148) );
  AOI22_X1 U74 ( .A1(DATA_OUT[16]), .A2(n94), .B1(DATA_IN[16]), .B2(n91), .ZN(
        n115) );
  INV_X1 U75 ( .A(n115), .ZN(n147) );
  AOI22_X1 U76 ( .A1(DATA_OUT[17]), .A2(n94), .B1(DATA_IN[17]), .B2(n91), .ZN(
        n116) );
  INV_X1 U77 ( .A(n116), .ZN(n146) );
  AOI22_X1 U78 ( .A1(DATA_OUT[18]), .A2(n94), .B1(DATA_IN[18]), .B2(n91), .ZN(
        n117) );
  INV_X1 U79 ( .A(n117), .ZN(n145) );
  AOI22_X1 U80 ( .A1(DATA_OUT[19]), .A2(n94), .B1(DATA_IN[19]), .B2(n91), .ZN(
        n118) );
  INV_X1 U81 ( .A(n118), .ZN(n144) );
  AOI22_X1 U82 ( .A1(DATA_OUT[20]), .A2(n94), .B1(DATA_IN[20]), .B2(n91), .ZN(
        n119) );
  INV_X1 U83 ( .A(n119), .ZN(n143) );
  AOI22_X1 U84 ( .A1(DATA_OUT[21]), .A2(n94), .B1(DATA_IN[21]), .B2(n91), .ZN(
        n120) );
  INV_X1 U85 ( .A(n120), .ZN(n142) );
  AOI22_X1 U86 ( .A1(DATA_OUT[22]), .A2(n94), .B1(DATA_IN[22]), .B2(n91), .ZN(
        n121) );
  INV_X1 U87 ( .A(n121), .ZN(n141) );
  AOI22_X1 U88 ( .A1(DATA_OUT[23]), .A2(n94), .B1(DATA_IN[23]), .B2(n91), .ZN(
        n122) );
  INV_X1 U89 ( .A(n122), .ZN(n140) );
  AOI22_X1 U90 ( .A1(DATA_OUT[24]), .A2(n95), .B1(DATA_IN[24]), .B2(n92), .ZN(
        n123) );
  INV_X1 U91 ( .A(n123), .ZN(n139) );
  AOI22_X1 U92 ( .A1(DATA_OUT[25]), .A2(n95), .B1(DATA_IN[25]), .B2(n92), .ZN(
        n124) );
  INV_X1 U93 ( .A(n124), .ZN(n138) );
  AOI22_X1 U94 ( .A1(DATA_OUT[26]), .A2(n95), .B1(DATA_IN[26]), .B2(n92), .ZN(
        n125) );
  INV_X1 U95 ( .A(n125), .ZN(n137) );
  AOI22_X1 U96 ( .A1(DATA_OUT[27]), .A2(n95), .B1(DATA_IN[27]), .B2(n92), .ZN(
        n126) );
  INV_X1 U97 ( .A(n126), .ZN(n136) );
  AOI22_X1 U98 ( .A1(DATA_OUT[28]), .A2(n95), .B1(DATA_IN[28]), .B2(n92), .ZN(
        n127) );
  INV_X1 U99 ( .A(n127), .ZN(n135) );
  AOI22_X1 U100 ( .A1(DATA_OUT[29]), .A2(n95), .B1(DATA_IN[29]), .B2(n92), 
        .ZN(n128) );
  INV_X1 U101 ( .A(n128), .ZN(n134) );
  AOI22_X1 U102 ( .A1(DATA_OUT[30]), .A2(n95), .B1(DATA_IN[30]), .B2(n92), 
        .ZN(n129) );
  INV_X1 U103 ( .A(n129), .ZN(n133) );
  AOI22_X1 U104 ( .A1(DATA_OUT[31]), .A2(n95), .B1(DATA_IN[31]), .B2(n92), 
        .ZN(n131) );
  INV_X1 U105 ( .A(n131), .ZN(n132) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n150), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n153), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n154), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n152), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n157), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n155), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n134), .CK(CLK), .Q(DATA_OUT[29]) );
  DFF_X1 \DATA_OUT_reg[28]  ( .D(n135), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X1 \DATA_OUT_reg[25]  ( .D(n138), .CK(CLK), .Q(DATA_OUT[25]) );
  DFF_X1 \DATA_OUT_reg[31]  ( .D(n132), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n133), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n137), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n139), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[23]  ( .D(n140), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n141), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n142), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n143), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n144), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n148), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n149), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n151), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n136), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n156), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n160), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n159), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n158), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n145), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n147), .CK(CLK), .Q(DATA_OUT[16]) );
endmodule


module REG_GENERIC_NBIT32_9 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;

  DFF_X1 \DATA_OUT_reg[31]  ( .D(n44), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n45), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n46), .CK(CLK), .Q(DATA_OUT[29]) );
  DFF_X1 \DATA_OUT_reg[28]  ( .D(n47), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n48), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n49), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[25]  ( .D(n50), .CK(CLK), .Q(DATA_OUT[25]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n51), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[23]  ( .D(n52), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n53), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n54), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n55), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n56), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n57), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n58), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n59), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n60), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n61), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n62), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n63), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n64), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n65), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n66), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n67), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n68), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n69), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n70), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n71), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n72), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n73), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n74), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n75), .CK(CLK), .Q(DATA_OUT[0]) );
  BUF_X2 U3 ( .A(n42), .Z(n5) );
  BUF_X2 U4 ( .A(n42), .Z(n6) );
  BUF_X1 U5 ( .A(n1), .Z(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n3) );
  BUF_X2 U7 ( .A(n42), .Z(n7) );
  BUF_X1 U8 ( .A(n1), .Z(n4) );
  AND2_X1 U9 ( .A1(n8), .A2(n10), .ZN(n1) );
  INV_X1 U10 ( .A(n9), .ZN(n8) );
  INV_X1 U11 ( .A(RST), .ZN(n9) );
  OR2_X1 U12 ( .A1(EN), .A2(n9), .ZN(n10) );
  INV_X1 U13 ( .A(n10), .ZN(n42) );
  AOI22_X1 U14 ( .A1(DATA_OUT[0]), .A2(n5), .B1(DATA_IN[0]), .B2(n2), .ZN(n11)
         );
  INV_X1 U15 ( .A(n11), .ZN(n75) );
  AOI22_X1 U16 ( .A1(DATA_OUT[1]), .A2(n5), .B1(DATA_IN[1]), .B2(n2), .ZN(n12)
         );
  INV_X1 U17 ( .A(n12), .ZN(n74) );
  AOI22_X1 U18 ( .A1(DATA_OUT[2]), .A2(n5), .B1(DATA_IN[2]), .B2(n2), .ZN(n13)
         );
  INV_X1 U19 ( .A(n13), .ZN(n73) );
  AOI22_X1 U20 ( .A1(DATA_OUT[3]), .A2(n5), .B1(DATA_IN[3]), .B2(n2), .ZN(n14)
         );
  INV_X1 U21 ( .A(n14), .ZN(n72) );
  AOI22_X1 U22 ( .A1(DATA_OUT[4]), .A2(n5), .B1(DATA_IN[4]), .B2(n2), .ZN(n15)
         );
  INV_X1 U23 ( .A(n15), .ZN(n71) );
  AOI22_X1 U24 ( .A1(DATA_OUT[5]), .A2(n5), .B1(DATA_IN[5]), .B2(n2), .ZN(n16)
         );
  INV_X1 U25 ( .A(n16), .ZN(n70) );
  AOI22_X1 U26 ( .A1(DATA_OUT[6]), .A2(n5), .B1(DATA_IN[6]), .B2(n2), .ZN(n17)
         );
  INV_X1 U27 ( .A(n17), .ZN(n69) );
  AOI22_X1 U28 ( .A1(DATA_OUT[7]), .A2(n5), .B1(DATA_IN[7]), .B2(n2), .ZN(n18)
         );
  INV_X1 U29 ( .A(n18), .ZN(n68) );
  AOI22_X1 U30 ( .A1(DATA_OUT[8]), .A2(n5), .B1(DATA_IN[8]), .B2(n2), .ZN(n19)
         );
  INV_X1 U31 ( .A(n19), .ZN(n67) );
  AOI22_X1 U32 ( .A1(DATA_OUT[9]), .A2(n5), .B1(DATA_IN[9]), .B2(n2), .ZN(n20)
         );
  INV_X1 U33 ( .A(n20), .ZN(n66) );
  AOI22_X1 U34 ( .A1(DATA_OUT[10]), .A2(n5), .B1(DATA_IN[10]), .B2(n2), .ZN(
        n21) );
  INV_X1 U35 ( .A(n21), .ZN(n65) );
  AOI22_X1 U36 ( .A1(DATA_OUT[11]), .A2(n5), .B1(DATA_IN[11]), .B2(n2), .ZN(
        n22) );
  INV_X1 U37 ( .A(n22), .ZN(n64) );
  AOI22_X1 U38 ( .A1(DATA_OUT[12]), .A2(n6), .B1(DATA_IN[12]), .B2(n3), .ZN(
        n23) );
  INV_X1 U39 ( .A(n23), .ZN(n63) );
  AOI22_X1 U40 ( .A1(DATA_OUT[13]), .A2(n6), .B1(DATA_IN[13]), .B2(n3), .ZN(
        n24) );
  INV_X1 U41 ( .A(n24), .ZN(n62) );
  AOI22_X1 U42 ( .A1(DATA_OUT[14]), .A2(n6), .B1(DATA_IN[14]), .B2(n3), .ZN(
        n25) );
  INV_X1 U43 ( .A(n25), .ZN(n61) );
  AOI22_X1 U44 ( .A1(DATA_OUT[15]), .A2(n6), .B1(DATA_IN[15]), .B2(n3), .ZN(
        n26) );
  INV_X1 U45 ( .A(n26), .ZN(n60) );
  AOI22_X1 U46 ( .A1(DATA_OUT[16]), .A2(n6), .B1(DATA_IN[16]), .B2(n3), .ZN(
        n27) );
  INV_X1 U47 ( .A(n27), .ZN(n59) );
  AOI22_X1 U48 ( .A1(DATA_OUT[17]), .A2(n6), .B1(DATA_IN[17]), .B2(n3), .ZN(
        n28) );
  INV_X1 U49 ( .A(n28), .ZN(n58) );
  AOI22_X1 U50 ( .A1(DATA_OUT[18]), .A2(n6), .B1(DATA_IN[18]), .B2(n3), .ZN(
        n29) );
  INV_X1 U51 ( .A(n29), .ZN(n57) );
  AOI22_X1 U52 ( .A1(DATA_OUT[19]), .A2(n6), .B1(DATA_IN[19]), .B2(n3), .ZN(
        n30) );
  INV_X1 U53 ( .A(n30), .ZN(n56) );
  AOI22_X1 U54 ( .A1(DATA_OUT[20]), .A2(n6), .B1(DATA_IN[20]), .B2(n3), .ZN(
        n31) );
  INV_X1 U55 ( .A(n31), .ZN(n55) );
  AOI22_X1 U56 ( .A1(DATA_OUT[21]), .A2(n6), .B1(DATA_IN[21]), .B2(n3), .ZN(
        n32) );
  INV_X1 U57 ( .A(n32), .ZN(n54) );
  AOI22_X1 U58 ( .A1(DATA_OUT[22]), .A2(n6), .B1(DATA_IN[22]), .B2(n3), .ZN(
        n33) );
  INV_X1 U59 ( .A(n33), .ZN(n53) );
  AOI22_X1 U60 ( .A1(DATA_OUT[23]), .A2(n6), .B1(DATA_IN[23]), .B2(n3), .ZN(
        n34) );
  INV_X1 U61 ( .A(n34), .ZN(n52) );
  AOI22_X1 U62 ( .A1(DATA_OUT[24]), .A2(n7), .B1(DATA_IN[24]), .B2(n4), .ZN(
        n35) );
  INV_X1 U63 ( .A(n35), .ZN(n51) );
  AOI22_X1 U64 ( .A1(DATA_OUT[25]), .A2(n7), .B1(DATA_IN[25]), .B2(n4), .ZN(
        n36) );
  INV_X1 U65 ( .A(n36), .ZN(n50) );
  AOI22_X1 U66 ( .A1(DATA_OUT[26]), .A2(n7), .B1(DATA_IN[26]), .B2(n4), .ZN(
        n37) );
  INV_X1 U67 ( .A(n37), .ZN(n49) );
  AOI22_X1 U68 ( .A1(DATA_OUT[27]), .A2(n7), .B1(DATA_IN[27]), .B2(n4), .ZN(
        n38) );
  INV_X1 U69 ( .A(n38), .ZN(n48) );
  AOI22_X1 U70 ( .A1(DATA_OUT[28]), .A2(n7), .B1(DATA_IN[28]), .B2(n4), .ZN(
        n39) );
  INV_X1 U71 ( .A(n39), .ZN(n47) );
  AOI22_X1 U72 ( .A1(DATA_OUT[29]), .A2(n7), .B1(DATA_IN[29]), .B2(n4), .ZN(
        n40) );
  INV_X1 U73 ( .A(n40), .ZN(n46) );
  AOI22_X1 U74 ( .A1(DATA_OUT[30]), .A2(n7), .B1(DATA_IN[30]), .B2(n4), .ZN(
        n41) );
  INV_X1 U75 ( .A(n41), .ZN(n45) );
  AOI22_X1 U76 ( .A1(DATA_OUT[31]), .A2(n7), .B1(DATA_IN[31]), .B2(n4), .ZN(
        n43) );
  INV_X1 U77 ( .A(n43), .ZN(n44) );
endmodule


module REG_GENERIC_NBIT32_8 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;

  DFF_X1 \DATA_OUT_reg[31]  ( .D(n44), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n45), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n46), .CK(CLK), .Q(DATA_OUT[29]) );
  DFF_X1 \DATA_OUT_reg[28]  ( .D(n47), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n48), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n49), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[25]  ( .D(n50), .CK(CLK), .Q(DATA_OUT[25]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n51), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[23]  ( .D(n52), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n53), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n54), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n55), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n56), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n57), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n58), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n59), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n60), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n61), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n62), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n63), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n64), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n65), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n66), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n67), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n68), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n69), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n70), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n71), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n72), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n73), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n74), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n75), .CK(CLK), .Q(DATA_OUT[0]) );
  BUF_X2 U3 ( .A(n42), .Z(n5) );
  BUF_X2 U4 ( .A(n42), .Z(n6) );
  BUF_X1 U5 ( .A(n1), .Z(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n3) );
  BUF_X2 U7 ( .A(n42), .Z(n7) );
  BUF_X1 U8 ( .A(n1), .Z(n4) );
  AND2_X1 U9 ( .A1(n8), .A2(n10), .ZN(n1) );
  INV_X1 U10 ( .A(n9), .ZN(n8) );
  INV_X1 U11 ( .A(RST), .ZN(n9) );
  OR2_X1 U12 ( .A1(EN), .A2(n9), .ZN(n10) );
  INV_X1 U13 ( .A(n10), .ZN(n42) );
  AOI22_X1 U14 ( .A1(DATA_OUT[0]), .A2(n5), .B1(DATA_IN[0]), .B2(n2), .ZN(n11)
         );
  INV_X1 U15 ( .A(n11), .ZN(n75) );
  AOI22_X1 U16 ( .A1(DATA_OUT[1]), .A2(n5), .B1(DATA_IN[1]), .B2(n2), .ZN(n12)
         );
  INV_X1 U17 ( .A(n12), .ZN(n74) );
  AOI22_X1 U18 ( .A1(DATA_OUT[2]), .A2(n5), .B1(DATA_IN[2]), .B2(n2), .ZN(n13)
         );
  INV_X1 U19 ( .A(n13), .ZN(n73) );
  AOI22_X1 U20 ( .A1(DATA_OUT[3]), .A2(n5), .B1(DATA_IN[3]), .B2(n2), .ZN(n14)
         );
  INV_X1 U21 ( .A(n14), .ZN(n72) );
  AOI22_X1 U22 ( .A1(DATA_OUT[4]), .A2(n5), .B1(DATA_IN[4]), .B2(n2), .ZN(n15)
         );
  INV_X1 U23 ( .A(n15), .ZN(n71) );
  AOI22_X1 U24 ( .A1(DATA_OUT[5]), .A2(n5), .B1(DATA_IN[5]), .B2(n2), .ZN(n16)
         );
  INV_X1 U25 ( .A(n16), .ZN(n70) );
  AOI22_X1 U26 ( .A1(DATA_OUT[6]), .A2(n5), .B1(DATA_IN[6]), .B2(n2), .ZN(n17)
         );
  INV_X1 U27 ( .A(n17), .ZN(n69) );
  AOI22_X1 U28 ( .A1(DATA_OUT[7]), .A2(n5), .B1(DATA_IN[7]), .B2(n2), .ZN(n18)
         );
  INV_X1 U29 ( .A(n18), .ZN(n68) );
  AOI22_X1 U30 ( .A1(DATA_OUT[8]), .A2(n5), .B1(DATA_IN[8]), .B2(n2), .ZN(n19)
         );
  INV_X1 U31 ( .A(n19), .ZN(n67) );
  AOI22_X1 U32 ( .A1(DATA_OUT[9]), .A2(n5), .B1(DATA_IN[9]), .B2(n2), .ZN(n20)
         );
  INV_X1 U33 ( .A(n20), .ZN(n66) );
  AOI22_X1 U34 ( .A1(DATA_OUT[10]), .A2(n5), .B1(DATA_IN[10]), .B2(n2), .ZN(
        n21) );
  INV_X1 U35 ( .A(n21), .ZN(n65) );
  AOI22_X1 U36 ( .A1(DATA_OUT[11]), .A2(n5), .B1(DATA_IN[11]), .B2(n2), .ZN(
        n22) );
  INV_X1 U37 ( .A(n22), .ZN(n64) );
  AOI22_X1 U38 ( .A1(DATA_OUT[12]), .A2(n6), .B1(DATA_IN[12]), .B2(n3), .ZN(
        n23) );
  INV_X1 U39 ( .A(n23), .ZN(n63) );
  AOI22_X1 U40 ( .A1(DATA_OUT[13]), .A2(n6), .B1(DATA_IN[13]), .B2(n3), .ZN(
        n24) );
  INV_X1 U41 ( .A(n24), .ZN(n62) );
  AOI22_X1 U42 ( .A1(DATA_OUT[14]), .A2(n6), .B1(DATA_IN[14]), .B2(n3), .ZN(
        n25) );
  INV_X1 U43 ( .A(n25), .ZN(n61) );
  AOI22_X1 U44 ( .A1(DATA_OUT[15]), .A2(n6), .B1(DATA_IN[15]), .B2(n3), .ZN(
        n26) );
  INV_X1 U45 ( .A(n26), .ZN(n60) );
  AOI22_X1 U46 ( .A1(DATA_OUT[16]), .A2(n6), .B1(DATA_IN[16]), .B2(n3), .ZN(
        n27) );
  INV_X1 U47 ( .A(n27), .ZN(n59) );
  AOI22_X1 U48 ( .A1(DATA_OUT[17]), .A2(n6), .B1(DATA_IN[17]), .B2(n3), .ZN(
        n28) );
  INV_X1 U49 ( .A(n28), .ZN(n58) );
  AOI22_X1 U50 ( .A1(DATA_OUT[18]), .A2(n6), .B1(DATA_IN[18]), .B2(n3), .ZN(
        n29) );
  INV_X1 U51 ( .A(n29), .ZN(n57) );
  AOI22_X1 U52 ( .A1(DATA_OUT[19]), .A2(n6), .B1(DATA_IN[19]), .B2(n3), .ZN(
        n30) );
  INV_X1 U53 ( .A(n30), .ZN(n56) );
  AOI22_X1 U54 ( .A1(DATA_OUT[20]), .A2(n6), .B1(DATA_IN[20]), .B2(n3), .ZN(
        n31) );
  INV_X1 U55 ( .A(n31), .ZN(n55) );
  AOI22_X1 U56 ( .A1(DATA_OUT[21]), .A2(n6), .B1(DATA_IN[21]), .B2(n3), .ZN(
        n32) );
  INV_X1 U57 ( .A(n32), .ZN(n54) );
  AOI22_X1 U58 ( .A1(DATA_OUT[22]), .A2(n6), .B1(DATA_IN[22]), .B2(n3), .ZN(
        n33) );
  INV_X1 U59 ( .A(n33), .ZN(n53) );
  AOI22_X1 U60 ( .A1(DATA_OUT[23]), .A2(n6), .B1(DATA_IN[23]), .B2(n3), .ZN(
        n34) );
  INV_X1 U61 ( .A(n34), .ZN(n52) );
  AOI22_X1 U62 ( .A1(DATA_OUT[24]), .A2(n7), .B1(DATA_IN[24]), .B2(n4), .ZN(
        n35) );
  INV_X1 U63 ( .A(n35), .ZN(n51) );
  AOI22_X1 U64 ( .A1(DATA_OUT[25]), .A2(n7), .B1(DATA_IN[25]), .B2(n4), .ZN(
        n36) );
  INV_X1 U65 ( .A(n36), .ZN(n50) );
  AOI22_X1 U66 ( .A1(DATA_OUT[26]), .A2(n7), .B1(DATA_IN[26]), .B2(n4), .ZN(
        n37) );
  INV_X1 U67 ( .A(n37), .ZN(n49) );
  AOI22_X1 U68 ( .A1(DATA_OUT[27]), .A2(n7), .B1(DATA_IN[27]), .B2(n4), .ZN(
        n38) );
  INV_X1 U69 ( .A(n38), .ZN(n48) );
  AOI22_X1 U70 ( .A1(DATA_OUT[28]), .A2(n7), .B1(DATA_IN[28]), .B2(n4), .ZN(
        n39) );
  INV_X1 U71 ( .A(n39), .ZN(n47) );
  AOI22_X1 U72 ( .A1(DATA_OUT[29]), .A2(n7), .B1(DATA_IN[29]), .B2(n4), .ZN(
        n40) );
  INV_X1 U73 ( .A(n40), .ZN(n46) );
  AOI22_X1 U74 ( .A1(DATA_OUT[30]), .A2(n7), .B1(DATA_IN[30]), .B2(n4), .ZN(
        n41) );
  INV_X1 U75 ( .A(n41), .ZN(n45) );
  AOI22_X1 U76 ( .A1(DATA_OUT[31]), .A2(n7), .B1(DATA_IN[31]), .B2(n4), .ZN(
        n43) );
  INV_X1 U77 ( .A(n43), .ZN(n44) );
endmodule


module REG_GENERIC_NBIT32_7 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;

  DFF_X1 \DATA_OUT_reg[31]  ( .D(n44), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n45), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n46), .CK(CLK), .Q(DATA_OUT[29]) );
  DFF_X1 \DATA_OUT_reg[28]  ( .D(n47), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n48), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n49), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[25]  ( .D(n50), .CK(CLK), .Q(DATA_OUT[25]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n51), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[23]  ( .D(n52), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n53), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n54), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n55), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n56), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n57), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n58), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n59), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n60), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n61), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n62), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n63), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n64), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n65), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n66), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n67), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n68), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n69), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n70), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n71), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n72), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n73), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n74), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n75), .CK(CLK), .Q(DATA_OUT[0]) );
  BUF_X2 U3 ( .A(n42), .Z(n5) );
  BUF_X2 U4 ( .A(n42), .Z(n6) );
  BUF_X1 U5 ( .A(n1), .Z(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n3) );
  BUF_X2 U7 ( .A(n42), .Z(n7) );
  BUF_X1 U8 ( .A(n1), .Z(n4) );
  AND2_X1 U9 ( .A1(n8), .A2(n10), .ZN(n1) );
  INV_X1 U10 ( .A(n9), .ZN(n8) );
  INV_X1 U11 ( .A(RST), .ZN(n9) );
  OR2_X1 U12 ( .A1(EN), .A2(n9), .ZN(n10) );
  INV_X1 U13 ( .A(n10), .ZN(n42) );
  AOI22_X1 U14 ( .A1(DATA_OUT[0]), .A2(n5), .B1(DATA_IN[0]), .B2(n2), .ZN(n11)
         );
  INV_X1 U15 ( .A(n11), .ZN(n75) );
  AOI22_X1 U16 ( .A1(DATA_OUT[1]), .A2(n5), .B1(DATA_IN[1]), .B2(n2), .ZN(n12)
         );
  INV_X1 U17 ( .A(n12), .ZN(n74) );
  AOI22_X1 U18 ( .A1(DATA_OUT[2]), .A2(n5), .B1(DATA_IN[2]), .B2(n2), .ZN(n13)
         );
  INV_X1 U19 ( .A(n13), .ZN(n73) );
  AOI22_X1 U20 ( .A1(DATA_OUT[3]), .A2(n5), .B1(DATA_IN[3]), .B2(n2), .ZN(n14)
         );
  INV_X1 U21 ( .A(n14), .ZN(n72) );
  AOI22_X1 U22 ( .A1(DATA_OUT[4]), .A2(n5), .B1(DATA_IN[4]), .B2(n2), .ZN(n15)
         );
  INV_X1 U23 ( .A(n15), .ZN(n71) );
  AOI22_X1 U24 ( .A1(DATA_OUT[5]), .A2(n5), .B1(DATA_IN[5]), .B2(n2), .ZN(n16)
         );
  INV_X1 U25 ( .A(n16), .ZN(n70) );
  AOI22_X1 U26 ( .A1(DATA_OUT[6]), .A2(n5), .B1(DATA_IN[6]), .B2(n2), .ZN(n17)
         );
  INV_X1 U27 ( .A(n17), .ZN(n69) );
  AOI22_X1 U28 ( .A1(DATA_OUT[7]), .A2(n5), .B1(DATA_IN[7]), .B2(n2), .ZN(n18)
         );
  INV_X1 U29 ( .A(n18), .ZN(n68) );
  AOI22_X1 U30 ( .A1(DATA_OUT[8]), .A2(n5), .B1(DATA_IN[8]), .B2(n2), .ZN(n19)
         );
  INV_X1 U31 ( .A(n19), .ZN(n67) );
  AOI22_X1 U32 ( .A1(DATA_OUT[9]), .A2(n5), .B1(DATA_IN[9]), .B2(n2), .ZN(n20)
         );
  INV_X1 U33 ( .A(n20), .ZN(n66) );
  AOI22_X1 U34 ( .A1(DATA_OUT[10]), .A2(n5), .B1(DATA_IN[10]), .B2(n2), .ZN(
        n21) );
  INV_X1 U35 ( .A(n21), .ZN(n65) );
  AOI22_X1 U36 ( .A1(DATA_OUT[11]), .A2(n5), .B1(DATA_IN[11]), .B2(n2), .ZN(
        n22) );
  INV_X1 U37 ( .A(n22), .ZN(n64) );
  AOI22_X1 U38 ( .A1(DATA_OUT[12]), .A2(n6), .B1(DATA_IN[12]), .B2(n3), .ZN(
        n23) );
  INV_X1 U39 ( .A(n23), .ZN(n63) );
  AOI22_X1 U40 ( .A1(DATA_OUT[13]), .A2(n6), .B1(DATA_IN[13]), .B2(n3), .ZN(
        n24) );
  INV_X1 U41 ( .A(n24), .ZN(n62) );
  AOI22_X1 U42 ( .A1(DATA_OUT[14]), .A2(n6), .B1(DATA_IN[14]), .B2(n3), .ZN(
        n25) );
  INV_X1 U43 ( .A(n25), .ZN(n61) );
  AOI22_X1 U44 ( .A1(DATA_OUT[15]), .A2(n6), .B1(DATA_IN[15]), .B2(n3), .ZN(
        n26) );
  INV_X1 U45 ( .A(n26), .ZN(n60) );
  AOI22_X1 U46 ( .A1(DATA_OUT[16]), .A2(n6), .B1(DATA_IN[16]), .B2(n3), .ZN(
        n27) );
  INV_X1 U47 ( .A(n27), .ZN(n59) );
  AOI22_X1 U48 ( .A1(DATA_OUT[17]), .A2(n6), .B1(DATA_IN[17]), .B2(n3), .ZN(
        n28) );
  INV_X1 U49 ( .A(n28), .ZN(n58) );
  AOI22_X1 U50 ( .A1(DATA_OUT[18]), .A2(n6), .B1(DATA_IN[18]), .B2(n3), .ZN(
        n29) );
  INV_X1 U51 ( .A(n29), .ZN(n57) );
  AOI22_X1 U52 ( .A1(DATA_OUT[19]), .A2(n6), .B1(DATA_IN[19]), .B2(n3), .ZN(
        n30) );
  INV_X1 U53 ( .A(n30), .ZN(n56) );
  AOI22_X1 U54 ( .A1(DATA_OUT[20]), .A2(n6), .B1(DATA_IN[20]), .B2(n3), .ZN(
        n31) );
  INV_X1 U55 ( .A(n31), .ZN(n55) );
  AOI22_X1 U56 ( .A1(DATA_OUT[21]), .A2(n6), .B1(DATA_IN[21]), .B2(n3), .ZN(
        n32) );
  INV_X1 U57 ( .A(n32), .ZN(n54) );
  AOI22_X1 U58 ( .A1(DATA_OUT[22]), .A2(n6), .B1(DATA_IN[22]), .B2(n3), .ZN(
        n33) );
  INV_X1 U59 ( .A(n33), .ZN(n53) );
  AOI22_X1 U60 ( .A1(DATA_OUT[23]), .A2(n6), .B1(DATA_IN[23]), .B2(n3), .ZN(
        n34) );
  INV_X1 U61 ( .A(n34), .ZN(n52) );
  AOI22_X1 U62 ( .A1(DATA_OUT[24]), .A2(n7), .B1(DATA_IN[24]), .B2(n4), .ZN(
        n35) );
  INV_X1 U63 ( .A(n35), .ZN(n51) );
  AOI22_X1 U64 ( .A1(DATA_OUT[25]), .A2(n7), .B1(DATA_IN[25]), .B2(n4), .ZN(
        n36) );
  INV_X1 U65 ( .A(n36), .ZN(n50) );
  AOI22_X1 U66 ( .A1(DATA_OUT[26]), .A2(n7), .B1(DATA_IN[26]), .B2(n4), .ZN(
        n37) );
  INV_X1 U67 ( .A(n37), .ZN(n49) );
  AOI22_X1 U68 ( .A1(DATA_OUT[27]), .A2(n7), .B1(DATA_IN[27]), .B2(n4), .ZN(
        n38) );
  INV_X1 U69 ( .A(n38), .ZN(n48) );
  AOI22_X1 U70 ( .A1(DATA_OUT[28]), .A2(n7), .B1(DATA_IN[28]), .B2(n4), .ZN(
        n39) );
  INV_X1 U71 ( .A(n39), .ZN(n47) );
  AOI22_X1 U72 ( .A1(DATA_OUT[29]), .A2(n7), .B1(DATA_IN[29]), .B2(n4), .ZN(
        n40) );
  INV_X1 U73 ( .A(n40), .ZN(n46) );
  AOI22_X1 U74 ( .A1(DATA_OUT[30]), .A2(n7), .B1(DATA_IN[30]), .B2(n4), .ZN(
        n41) );
  INV_X1 U75 ( .A(n41), .ZN(n45) );
  AOI22_X1 U76 ( .A1(DATA_OUT[31]), .A2(n7), .B1(DATA_IN[31]), .B2(n4), .ZN(
        n43) );
  INV_X1 U77 ( .A(n43), .ZN(n44) );
endmodule


module REG_GENERIC_NBIT32_6 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;

  DFF_X1 \DATA_OUT_reg[31]  ( .D(n44), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n45), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n46), .CK(CLK), .Q(DATA_OUT[29]) );
  DFF_X1 \DATA_OUT_reg[28]  ( .D(n47), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n48), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n49), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[25]  ( .D(n50), .CK(CLK), .Q(DATA_OUT[25]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n51), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[23]  ( .D(n52), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n53), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n54), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n55), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n56), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n57), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n58), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n59), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n60), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n61), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n62), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n63), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n64), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n65), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n66), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n67), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n68), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n69), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n70), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n71), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n72), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n73), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n74), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n75), .CK(CLK), .Q(DATA_OUT[0]) );
  BUF_X2 U3 ( .A(n42), .Z(n5) );
  BUF_X2 U4 ( .A(n42), .Z(n6) );
  BUF_X1 U5 ( .A(n1), .Z(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n3) );
  BUF_X2 U7 ( .A(n42), .Z(n7) );
  BUF_X1 U8 ( .A(n1), .Z(n4) );
  AND2_X1 U9 ( .A1(n8), .A2(n10), .ZN(n1) );
  INV_X1 U10 ( .A(n9), .ZN(n8) );
  INV_X1 U11 ( .A(RST), .ZN(n9) );
  OR2_X1 U12 ( .A1(EN), .A2(n9), .ZN(n10) );
  INV_X1 U13 ( .A(n10), .ZN(n42) );
  AOI22_X1 U14 ( .A1(DATA_OUT[0]), .A2(n5), .B1(DATA_IN[0]), .B2(n2), .ZN(n11)
         );
  INV_X1 U15 ( .A(n11), .ZN(n75) );
  AOI22_X1 U16 ( .A1(DATA_OUT[1]), .A2(n5), .B1(DATA_IN[1]), .B2(n2), .ZN(n12)
         );
  INV_X1 U17 ( .A(n12), .ZN(n74) );
  AOI22_X1 U18 ( .A1(DATA_OUT[2]), .A2(n5), .B1(DATA_IN[2]), .B2(n2), .ZN(n13)
         );
  INV_X1 U19 ( .A(n13), .ZN(n73) );
  AOI22_X1 U20 ( .A1(DATA_OUT[3]), .A2(n5), .B1(DATA_IN[3]), .B2(n2), .ZN(n14)
         );
  INV_X1 U21 ( .A(n14), .ZN(n72) );
  AOI22_X1 U22 ( .A1(DATA_OUT[4]), .A2(n5), .B1(DATA_IN[4]), .B2(n2), .ZN(n15)
         );
  INV_X1 U23 ( .A(n15), .ZN(n71) );
  AOI22_X1 U24 ( .A1(DATA_OUT[5]), .A2(n5), .B1(DATA_IN[5]), .B2(n2), .ZN(n16)
         );
  INV_X1 U25 ( .A(n16), .ZN(n70) );
  AOI22_X1 U26 ( .A1(DATA_OUT[6]), .A2(n5), .B1(DATA_IN[6]), .B2(n2), .ZN(n17)
         );
  INV_X1 U27 ( .A(n17), .ZN(n69) );
  AOI22_X1 U28 ( .A1(DATA_OUT[7]), .A2(n5), .B1(DATA_IN[7]), .B2(n2), .ZN(n18)
         );
  INV_X1 U29 ( .A(n18), .ZN(n68) );
  AOI22_X1 U30 ( .A1(DATA_OUT[8]), .A2(n5), .B1(DATA_IN[8]), .B2(n2), .ZN(n19)
         );
  INV_X1 U31 ( .A(n19), .ZN(n67) );
  AOI22_X1 U32 ( .A1(DATA_OUT[9]), .A2(n5), .B1(DATA_IN[9]), .B2(n2), .ZN(n20)
         );
  INV_X1 U33 ( .A(n20), .ZN(n66) );
  AOI22_X1 U34 ( .A1(DATA_OUT[10]), .A2(n5), .B1(DATA_IN[10]), .B2(n2), .ZN(
        n21) );
  INV_X1 U35 ( .A(n21), .ZN(n65) );
  AOI22_X1 U36 ( .A1(DATA_OUT[11]), .A2(n5), .B1(DATA_IN[11]), .B2(n2), .ZN(
        n22) );
  INV_X1 U37 ( .A(n22), .ZN(n64) );
  AOI22_X1 U38 ( .A1(DATA_OUT[12]), .A2(n6), .B1(DATA_IN[12]), .B2(n3), .ZN(
        n23) );
  INV_X1 U39 ( .A(n23), .ZN(n63) );
  AOI22_X1 U40 ( .A1(DATA_OUT[13]), .A2(n6), .B1(DATA_IN[13]), .B2(n3), .ZN(
        n24) );
  INV_X1 U41 ( .A(n24), .ZN(n62) );
  AOI22_X1 U42 ( .A1(DATA_OUT[14]), .A2(n6), .B1(DATA_IN[14]), .B2(n3), .ZN(
        n25) );
  INV_X1 U43 ( .A(n25), .ZN(n61) );
  AOI22_X1 U44 ( .A1(DATA_OUT[15]), .A2(n6), .B1(DATA_IN[15]), .B2(n3), .ZN(
        n26) );
  INV_X1 U45 ( .A(n26), .ZN(n60) );
  AOI22_X1 U46 ( .A1(DATA_OUT[16]), .A2(n6), .B1(DATA_IN[16]), .B2(n3), .ZN(
        n27) );
  INV_X1 U47 ( .A(n27), .ZN(n59) );
  AOI22_X1 U48 ( .A1(DATA_OUT[17]), .A2(n6), .B1(DATA_IN[17]), .B2(n3), .ZN(
        n28) );
  INV_X1 U49 ( .A(n28), .ZN(n58) );
  AOI22_X1 U50 ( .A1(DATA_OUT[18]), .A2(n6), .B1(DATA_IN[18]), .B2(n3), .ZN(
        n29) );
  INV_X1 U51 ( .A(n29), .ZN(n57) );
  AOI22_X1 U52 ( .A1(DATA_OUT[19]), .A2(n6), .B1(DATA_IN[19]), .B2(n3), .ZN(
        n30) );
  INV_X1 U53 ( .A(n30), .ZN(n56) );
  AOI22_X1 U54 ( .A1(DATA_OUT[20]), .A2(n6), .B1(DATA_IN[20]), .B2(n3), .ZN(
        n31) );
  INV_X1 U55 ( .A(n31), .ZN(n55) );
  AOI22_X1 U56 ( .A1(DATA_OUT[21]), .A2(n6), .B1(DATA_IN[21]), .B2(n3), .ZN(
        n32) );
  INV_X1 U57 ( .A(n32), .ZN(n54) );
  AOI22_X1 U58 ( .A1(DATA_OUT[22]), .A2(n6), .B1(DATA_IN[22]), .B2(n3), .ZN(
        n33) );
  INV_X1 U59 ( .A(n33), .ZN(n53) );
  AOI22_X1 U60 ( .A1(DATA_OUT[23]), .A2(n6), .B1(DATA_IN[23]), .B2(n3), .ZN(
        n34) );
  INV_X1 U61 ( .A(n34), .ZN(n52) );
  AOI22_X1 U62 ( .A1(DATA_OUT[24]), .A2(n7), .B1(DATA_IN[24]), .B2(n4), .ZN(
        n35) );
  INV_X1 U63 ( .A(n35), .ZN(n51) );
  AOI22_X1 U64 ( .A1(DATA_OUT[25]), .A2(n7), .B1(DATA_IN[25]), .B2(n4), .ZN(
        n36) );
  INV_X1 U65 ( .A(n36), .ZN(n50) );
  AOI22_X1 U66 ( .A1(DATA_OUT[26]), .A2(n7), .B1(DATA_IN[26]), .B2(n4), .ZN(
        n37) );
  INV_X1 U67 ( .A(n37), .ZN(n49) );
  AOI22_X1 U68 ( .A1(DATA_OUT[27]), .A2(n7), .B1(DATA_IN[27]), .B2(n4), .ZN(
        n38) );
  INV_X1 U69 ( .A(n38), .ZN(n48) );
  AOI22_X1 U70 ( .A1(DATA_OUT[28]), .A2(n7), .B1(DATA_IN[28]), .B2(n4), .ZN(
        n39) );
  INV_X1 U71 ( .A(n39), .ZN(n47) );
  AOI22_X1 U72 ( .A1(DATA_OUT[29]), .A2(n7), .B1(DATA_IN[29]), .B2(n4), .ZN(
        n40) );
  INV_X1 U73 ( .A(n40), .ZN(n46) );
  AOI22_X1 U74 ( .A1(DATA_OUT[30]), .A2(n7), .B1(DATA_IN[30]), .B2(n4), .ZN(
        n41) );
  INV_X1 U75 ( .A(n41), .ZN(n45) );
  AOI22_X1 U76 ( .A1(DATA_OUT[31]), .A2(n7), .B1(DATA_IN[31]), .B2(n4), .ZN(
        n43) );
  INV_X1 U77 ( .A(n43), .ZN(n44) );
endmodule


module REG_GENERIC_NBIT32_5 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;

  DFF_X1 \DATA_OUT_reg[31]  ( .D(n44), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n45), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n48), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n49), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n51), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n53), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n54), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n55), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n56), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n57), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n58), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n59), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n60), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n61), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n62), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n63), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n64), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n65), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n66), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n67), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n68), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n69), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n70), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n71), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n72), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n73), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n74), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n75), .CK(CLK), .Q(DATA_OUT[0]) );
  DFF_X2 \DATA_OUT_reg[23]  ( .D(n52), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X2 \DATA_OUT_reg[28]  ( .D(n47), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X2 \DATA_OUT_reg[25]  ( .D(n50), .CK(CLK), .Q(DATA_OUT[25]) );
  BUF_X2 U3 ( .A(n42), .Z(n5) );
  BUF_X2 U4 ( .A(n42), .Z(n6) );
  BUF_X1 U5 ( .A(n1), .Z(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n3) );
  BUF_X2 U7 ( .A(n42), .Z(n7) );
  BUF_X1 U8 ( .A(n1), .Z(n4) );
  AND2_X1 U9 ( .A1(n8), .A2(n10), .ZN(n1) );
  INV_X1 U10 ( .A(n9), .ZN(n8) );
  INV_X1 U11 ( .A(RST), .ZN(n9) );
  OR2_X1 U12 ( .A1(EN), .A2(n9), .ZN(n10) );
  INV_X1 U13 ( .A(n10), .ZN(n42) );
  AOI22_X1 U14 ( .A1(DATA_OUT[0]), .A2(n5), .B1(DATA_IN[0]), .B2(n2), .ZN(n11)
         );
  INV_X1 U15 ( .A(n11), .ZN(n75) );
  AOI22_X1 U16 ( .A1(DATA_OUT[1]), .A2(n5), .B1(DATA_IN[1]), .B2(n2), .ZN(n12)
         );
  INV_X1 U17 ( .A(n12), .ZN(n74) );
  AOI22_X1 U18 ( .A1(DATA_OUT[2]), .A2(n5), .B1(DATA_IN[2]), .B2(n2), .ZN(n13)
         );
  INV_X1 U19 ( .A(n13), .ZN(n73) );
  AOI22_X1 U20 ( .A1(DATA_OUT[3]), .A2(n5), .B1(DATA_IN[3]), .B2(n2), .ZN(n14)
         );
  INV_X1 U21 ( .A(n14), .ZN(n72) );
  AOI22_X1 U22 ( .A1(DATA_OUT[4]), .A2(n5), .B1(DATA_IN[4]), .B2(n2), .ZN(n15)
         );
  INV_X1 U23 ( .A(n15), .ZN(n71) );
  AOI22_X1 U24 ( .A1(DATA_OUT[5]), .A2(n5), .B1(DATA_IN[5]), .B2(n2), .ZN(n16)
         );
  INV_X1 U25 ( .A(n16), .ZN(n70) );
  AOI22_X1 U26 ( .A1(DATA_OUT[6]), .A2(n5), .B1(DATA_IN[6]), .B2(n2), .ZN(n17)
         );
  INV_X1 U27 ( .A(n17), .ZN(n69) );
  AOI22_X1 U28 ( .A1(DATA_OUT[7]), .A2(n5), .B1(DATA_IN[7]), .B2(n2), .ZN(n18)
         );
  INV_X1 U29 ( .A(n18), .ZN(n68) );
  AOI22_X1 U30 ( .A1(DATA_OUT[8]), .A2(n5), .B1(DATA_IN[8]), .B2(n2), .ZN(n19)
         );
  INV_X1 U31 ( .A(n19), .ZN(n67) );
  AOI22_X1 U32 ( .A1(DATA_OUT[9]), .A2(n5), .B1(DATA_IN[9]), .B2(n2), .ZN(n20)
         );
  INV_X1 U33 ( .A(n20), .ZN(n66) );
  AOI22_X1 U34 ( .A1(DATA_OUT[10]), .A2(n5), .B1(DATA_IN[10]), .B2(n2), .ZN(
        n21) );
  INV_X1 U35 ( .A(n21), .ZN(n65) );
  AOI22_X1 U36 ( .A1(DATA_OUT[11]), .A2(n5), .B1(DATA_IN[11]), .B2(n2), .ZN(
        n22) );
  INV_X1 U37 ( .A(n22), .ZN(n64) );
  AOI22_X1 U38 ( .A1(DATA_OUT[12]), .A2(n6), .B1(DATA_IN[12]), .B2(n3), .ZN(
        n23) );
  INV_X1 U39 ( .A(n23), .ZN(n63) );
  AOI22_X1 U40 ( .A1(DATA_OUT[13]), .A2(n6), .B1(DATA_IN[13]), .B2(n3), .ZN(
        n24) );
  INV_X1 U41 ( .A(n24), .ZN(n62) );
  AOI22_X1 U42 ( .A1(DATA_OUT[14]), .A2(n6), .B1(DATA_IN[14]), .B2(n3), .ZN(
        n25) );
  INV_X1 U43 ( .A(n25), .ZN(n61) );
  AOI22_X1 U44 ( .A1(DATA_OUT[15]), .A2(n6), .B1(DATA_IN[15]), .B2(n3), .ZN(
        n26) );
  INV_X1 U45 ( .A(n26), .ZN(n60) );
  AOI22_X1 U46 ( .A1(DATA_OUT[16]), .A2(n6), .B1(DATA_IN[16]), .B2(n3), .ZN(
        n27) );
  INV_X1 U47 ( .A(n27), .ZN(n59) );
  AOI22_X1 U48 ( .A1(DATA_OUT[17]), .A2(n6), .B1(DATA_IN[17]), .B2(n3), .ZN(
        n28) );
  INV_X1 U49 ( .A(n28), .ZN(n58) );
  AOI22_X1 U50 ( .A1(DATA_OUT[18]), .A2(n6), .B1(DATA_IN[18]), .B2(n3), .ZN(
        n29) );
  INV_X1 U51 ( .A(n29), .ZN(n57) );
  AOI22_X1 U52 ( .A1(DATA_OUT[19]), .A2(n6), .B1(DATA_IN[19]), .B2(n3), .ZN(
        n30) );
  INV_X1 U53 ( .A(n30), .ZN(n56) );
  AOI22_X1 U54 ( .A1(DATA_OUT[20]), .A2(n6), .B1(DATA_IN[20]), .B2(n3), .ZN(
        n31) );
  INV_X1 U55 ( .A(n31), .ZN(n55) );
  AOI22_X1 U56 ( .A1(DATA_OUT[21]), .A2(n6), .B1(DATA_IN[21]), .B2(n3), .ZN(
        n32) );
  INV_X1 U57 ( .A(n32), .ZN(n54) );
  AOI22_X1 U58 ( .A1(DATA_OUT[22]), .A2(n6), .B1(DATA_IN[22]), .B2(n3), .ZN(
        n33) );
  INV_X1 U59 ( .A(n33), .ZN(n53) );
  AOI22_X1 U60 ( .A1(DATA_OUT[23]), .A2(n6), .B1(DATA_IN[23]), .B2(n3), .ZN(
        n34) );
  INV_X1 U61 ( .A(n34), .ZN(n52) );
  AOI22_X1 U62 ( .A1(DATA_OUT[24]), .A2(n7), .B1(DATA_IN[24]), .B2(n4), .ZN(
        n35) );
  INV_X1 U63 ( .A(n35), .ZN(n51) );
  AOI22_X1 U64 ( .A1(DATA_OUT[25]), .A2(n7), .B1(DATA_IN[25]), .B2(n4), .ZN(
        n36) );
  INV_X1 U65 ( .A(n36), .ZN(n50) );
  AOI22_X1 U66 ( .A1(DATA_OUT[26]), .A2(n7), .B1(DATA_IN[26]), .B2(n4), .ZN(
        n37) );
  INV_X1 U67 ( .A(n37), .ZN(n49) );
  AOI22_X1 U68 ( .A1(DATA_OUT[27]), .A2(n7), .B1(DATA_IN[27]), .B2(n4), .ZN(
        n38) );
  INV_X1 U69 ( .A(n38), .ZN(n48) );
  AOI22_X1 U70 ( .A1(DATA_OUT[28]), .A2(n7), .B1(DATA_IN[28]), .B2(n4), .ZN(
        n39) );
  INV_X1 U71 ( .A(n39), .ZN(n47) );
  AOI22_X1 U72 ( .A1(DATA_OUT[29]), .A2(n7), .B1(DATA_IN[29]), .B2(n4), .ZN(
        n40) );
  INV_X1 U73 ( .A(n40), .ZN(n46) );
  AOI22_X1 U74 ( .A1(DATA_OUT[30]), .A2(n7), .B1(DATA_IN[30]), .B2(n4), .ZN(
        n41) );
  INV_X1 U75 ( .A(n41), .ZN(n45) );
  AOI22_X1 U76 ( .A1(DATA_OUT[31]), .A2(n7), .B1(DATA_IN[31]), .B2(n4), .ZN(
        n43) );
  INV_X1 U77 ( .A(n43), .ZN(n44) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n46), .CK(CLK), .Q(DATA_OUT[29]) );
endmodule


module REG_GENERIC_NBIT32_4 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;

  DFF_X1 \DATA_OUT_reg[31]  ( .D(n44), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n45), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n46), .CK(CLK), .Q(DATA_OUT[29]) );
  DFF_X1 \DATA_OUT_reg[28]  ( .D(n47), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n48), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n49), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[25]  ( .D(n50), .CK(CLK), .Q(DATA_OUT[25]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n51), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[23]  ( .D(n52), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n53), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n54), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n55), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n56), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n57), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n58), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n59), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n60), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n61), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n62), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n63), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n64), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n65), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n66), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n67), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n68), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n69), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n70), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n71), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n72), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n73), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n74), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n75), .CK(CLK), .Q(DATA_OUT[0]) );
  BUF_X2 U3 ( .A(n42), .Z(n6) );
  BUF_X2 U4 ( .A(n42), .Z(n5) );
  BUF_X1 U5 ( .A(n1), .Z(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n3) );
  BUF_X2 U7 ( .A(n42), .Z(n7) );
  BUF_X1 U8 ( .A(n1), .Z(n4) );
  AND2_X1 U9 ( .A1(n8), .A2(n10), .ZN(n1) );
  INV_X1 U10 ( .A(n9), .ZN(n8) );
  INV_X1 U11 ( .A(RST), .ZN(n9) );
  OR2_X1 U12 ( .A1(EN), .A2(n9), .ZN(n10) );
  INV_X1 U13 ( .A(n10), .ZN(n42) );
  AOI22_X1 U14 ( .A1(DATA_OUT[0]), .A2(n5), .B1(DATA_IN[0]), .B2(n2), .ZN(n11)
         );
  INV_X1 U15 ( .A(n11), .ZN(n75) );
  AOI22_X1 U16 ( .A1(DATA_OUT[1]), .A2(n5), .B1(DATA_IN[1]), .B2(n2), .ZN(n12)
         );
  INV_X1 U17 ( .A(n12), .ZN(n74) );
  AOI22_X1 U18 ( .A1(DATA_OUT[2]), .A2(n5), .B1(DATA_IN[2]), .B2(n2), .ZN(n13)
         );
  INV_X1 U19 ( .A(n13), .ZN(n73) );
  AOI22_X1 U20 ( .A1(DATA_OUT[3]), .A2(n5), .B1(DATA_IN[3]), .B2(n2), .ZN(n14)
         );
  INV_X1 U21 ( .A(n14), .ZN(n72) );
  AOI22_X1 U22 ( .A1(DATA_OUT[4]), .A2(n5), .B1(DATA_IN[4]), .B2(n2), .ZN(n15)
         );
  INV_X1 U23 ( .A(n15), .ZN(n71) );
  AOI22_X1 U24 ( .A1(DATA_OUT[5]), .A2(n5), .B1(DATA_IN[5]), .B2(n2), .ZN(n16)
         );
  INV_X1 U25 ( .A(n16), .ZN(n70) );
  AOI22_X1 U26 ( .A1(DATA_OUT[6]), .A2(n5), .B1(DATA_IN[6]), .B2(n2), .ZN(n17)
         );
  INV_X1 U27 ( .A(n17), .ZN(n69) );
  AOI22_X1 U28 ( .A1(DATA_OUT[7]), .A2(n5), .B1(DATA_IN[7]), .B2(n2), .ZN(n18)
         );
  INV_X1 U29 ( .A(n18), .ZN(n68) );
  AOI22_X1 U30 ( .A1(DATA_OUT[8]), .A2(n5), .B1(DATA_IN[8]), .B2(n2), .ZN(n19)
         );
  INV_X1 U31 ( .A(n19), .ZN(n67) );
  AOI22_X1 U32 ( .A1(DATA_OUT[9]), .A2(n5), .B1(DATA_IN[9]), .B2(n2), .ZN(n20)
         );
  INV_X1 U33 ( .A(n20), .ZN(n66) );
  AOI22_X1 U34 ( .A1(DATA_OUT[10]), .A2(n5), .B1(DATA_IN[10]), .B2(n2), .ZN(
        n21) );
  INV_X1 U35 ( .A(n21), .ZN(n65) );
  AOI22_X1 U36 ( .A1(DATA_OUT[11]), .A2(n5), .B1(DATA_IN[11]), .B2(n2), .ZN(
        n22) );
  INV_X1 U37 ( .A(n22), .ZN(n64) );
  AOI22_X1 U38 ( .A1(DATA_OUT[12]), .A2(n6), .B1(DATA_IN[12]), .B2(n3), .ZN(
        n23) );
  INV_X1 U39 ( .A(n23), .ZN(n63) );
  AOI22_X1 U40 ( .A1(DATA_OUT[13]), .A2(n6), .B1(DATA_IN[13]), .B2(n3), .ZN(
        n24) );
  INV_X1 U41 ( .A(n24), .ZN(n62) );
  AOI22_X1 U42 ( .A1(DATA_OUT[14]), .A2(n6), .B1(DATA_IN[14]), .B2(n3), .ZN(
        n25) );
  INV_X1 U43 ( .A(n25), .ZN(n61) );
  AOI22_X1 U44 ( .A1(DATA_OUT[15]), .A2(n6), .B1(DATA_IN[15]), .B2(n3), .ZN(
        n26) );
  INV_X1 U45 ( .A(n26), .ZN(n60) );
  AOI22_X1 U46 ( .A1(DATA_OUT[16]), .A2(n6), .B1(DATA_IN[16]), .B2(n3), .ZN(
        n27) );
  INV_X1 U47 ( .A(n27), .ZN(n59) );
  AOI22_X1 U48 ( .A1(DATA_OUT[17]), .A2(n6), .B1(DATA_IN[17]), .B2(n3), .ZN(
        n28) );
  INV_X1 U49 ( .A(n28), .ZN(n58) );
  AOI22_X1 U50 ( .A1(DATA_OUT[18]), .A2(n6), .B1(DATA_IN[18]), .B2(n3), .ZN(
        n29) );
  INV_X1 U51 ( .A(n29), .ZN(n57) );
  AOI22_X1 U52 ( .A1(DATA_OUT[19]), .A2(n6), .B1(DATA_IN[19]), .B2(n3), .ZN(
        n30) );
  INV_X1 U53 ( .A(n30), .ZN(n56) );
  AOI22_X1 U54 ( .A1(DATA_OUT[20]), .A2(n6), .B1(DATA_IN[20]), .B2(n3), .ZN(
        n31) );
  INV_X1 U55 ( .A(n31), .ZN(n55) );
  AOI22_X1 U56 ( .A1(DATA_OUT[21]), .A2(n6), .B1(DATA_IN[21]), .B2(n3), .ZN(
        n32) );
  INV_X1 U57 ( .A(n32), .ZN(n54) );
  AOI22_X1 U58 ( .A1(DATA_OUT[22]), .A2(n6), .B1(DATA_IN[22]), .B2(n3), .ZN(
        n33) );
  INV_X1 U59 ( .A(n33), .ZN(n53) );
  AOI22_X1 U60 ( .A1(DATA_OUT[23]), .A2(n6), .B1(DATA_IN[23]), .B2(n3), .ZN(
        n34) );
  INV_X1 U61 ( .A(n34), .ZN(n52) );
  AOI22_X1 U62 ( .A1(DATA_OUT[24]), .A2(n7), .B1(DATA_IN[24]), .B2(n4), .ZN(
        n35) );
  INV_X1 U63 ( .A(n35), .ZN(n51) );
  AOI22_X1 U64 ( .A1(DATA_OUT[25]), .A2(n7), .B1(DATA_IN[25]), .B2(n4), .ZN(
        n36) );
  INV_X1 U65 ( .A(n36), .ZN(n50) );
  AOI22_X1 U66 ( .A1(DATA_OUT[26]), .A2(n7), .B1(DATA_IN[26]), .B2(n4), .ZN(
        n37) );
  INV_X1 U67 ( .A(n37), .ZN(n49) );
  AOI22_X1 U68 ( .A1(DATA_OUT[27]), .A2(n7), .B1(DATA_IN[27]), .B2(n4), .ZN(
        n38) );
  INV_X1 U69 ( .A(n38), .ZN(n48) );
  AOI22_X1 U70 ( .A1(DATA_OUT[28]), .A2(n7), .B1(DATA_IN[28]), .B2(n4), .ZN(
        n39) );
  INV_X1 U71 ( .A(n39), .ZN(n47) );
  AOI22_X1 U72 ( .A1(DATA_OUT[29]), .A2(n7), .B1(DATA_IN[29]), .B2(n4), .ZN(
        n40) );
  INV_X1 U73 ( .A(n40), .ZN(n46) );
  AOI22_X1 U74 ( .A1(DATA_OUT[30]), .A2(n7), .B1(DATA_IN[30]), .B2(n4), .ZN(
        n41) );
  INV_X1 U75 ( .A(n41), .ZN(n45) );
  AOI22_X1 U76 ( .A1(DATA_OUT[31]), .A2(n7), .B1(DATA_IN[31]), .B2(n4), .ZN(
        n43) );
  INV_X1 U77 ( .A(n43), .ZN(n44) );
endmodule


module REG_GENERIC_NBIT26 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [25:0] DATA_IN;
  output [25:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;

  DFF_X1 \DATA_OUT_reg[25]  ( .D(n38), .CK(CLK), .Q(DATA_OUT[25]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n39), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[23]  ( .D(n40), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n41), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n42), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n43), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n44), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n45), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n46), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n47), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n48), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n49), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n50), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n51), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n52), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n53), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n54), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n55), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n56), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n57), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n58), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n59), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n60), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n61), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n62), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n63), .CK(CLK), .Q(DATA_OUT[0]) );
  CLKBUF_X1 U3 ( .A(n1), .Z(n4) );
  BUF_X1 U4 ( .A(n36), .Z(n5) );
  BUF_X1 U5 ( .A(n36), .Z(n6) );
  BUF_X1 U6 ( .A(n1), .Z(n3) );
  BUF_X1 U7 ( .A(n1), .Z(n2) );
  CLKBUF_X1 U8 ( .A(n36), .Z(n7) );
  AND2_X1 U9 ( .A1(n8), .A2(n10), .ZN(n1) );
  INV_X1 U10 ( .A(n9), .ZN(n8) );
  INV_X1 U11 ( .A(RST), .ZN(n9) );
  OR2_X1 U12 ( .A1(EN), .A2(n9), .ZN(n10) );
  INV_X1 U13 ( .A(n10), .ZN(n36) );
  AOI22_X1 U14 ( .A1(DATA_OUT[0]), .A2(n5), .B1(DATA_IN[0]), .B2(n4), .ZN(n11)
         );
  INV_X1 U15 ( .A(n11), .ZN(n63) );
  AOI22_X1 U16 ( .A1(DATA_OUT[1]), .A2(n5), .B1(DATA_IN[1]), .B2(n4), .ZN(n12)
         );
  INV_X1 U17 ( .A(n12), .ZN(n62) );
  AOI22_X1 U18 ( .A1(DATA_OUT[2]), .A2(n5), .B1(DATA_IN[2]), .B2(n3), .ZN(n13)
         );
  INV_X1 U19 ( .A(n13), .ZN(n61) );
  AOI22_X1 U20 ( .A1(DATA_OUT[3]), .A2(n5), .B1(DATA_IN[3]), .B2(n3), .ZN(n14)
         );
  INV_X1 U21 ( .A(n14), .ZN(n60) );
  AOI22_X1 U22 ( .A1(DATA_OUT[4]), .A2(n5), .B1(DATA_IN[4]), .B2(n3), .ZN(n15)
         );
  INV_X1 U23 ( .A(n15), .ZN(n59) );
  AOI22_X1 U24 ( .A1(DATA_OUT[5]), .A2(n5), .B1(DATA_IN[5]), .B2(n3), .ZN(n16)
         );
  INV_X1 U25 ( .A(n16), .ZN(n58) );
  AOI22_X1 U26 ( .A1(DATA_OUT[6]), .A2(n5), .B1(DATA_IN[6]), .B2(n3), .ZN(n17)
         );
  INV_X1 U27 ( .A(n17), .ZN(n57) );
  AOI22_X1 U28 ( .A1(DATA_OUT[7]), .A2(n5), .B1(DATA_IN[7]), .B2(n3), .ZN(n18)
         );
  INV_X1 U29 ( .A(n18), .ZN(n56) );
  AOI22_X1 U30 ( .A1(DATA_OUT[8]), .A2(n5), .B1(DATA_IN[8]), .B2(n3), .ZN(n19)
         );
  INV_X1 U31 ( .A(n19), .ZN(n55) );
  AOI22_X1 U32 ( .A1(DATA_OUT[9]), .A2(n5), .B1(DATA_IN[9]), .B2(n3), .ZN(n20)
         );
  INV_X1 U33 ( .A(n20), .ZN(n54) );
  AOI22_X1 U34 ( .A1(DATA_OUT[10]), .A2(n5), .B1(DATA_IN[10]), .B2(n3), .ZN(
        n21) );
  INV_X1 U35 ( .A(n21), .ZN(n53) );
  AOI22_X1 U36 ( .A1(DATA_OUT[11]), .A2(n5), .B1(DATA_IN[11]), .B2(n3), .ZN(
        n22) );
  INV_X1 U37 ( .A(n22), .ZN(n52) );
  AOI22_X1 U38 ( .A1(DATA_OUT[12]), .A2(n6), .B1(DATA_IN[12]), .B2(n3), .ZN(
        n23) );
  INV_X1 U39 ( .A(n23), .ZN(n51) );
  AOI22_X1 U40 ( .A1(DATA_OUT[13]), .A2(n6), .B1(DATA_IN[13]), .B2(n3), .ZN(
        n24) );
  INV_X1 U41 ( .A(n24), .ZN(n50) );
  AOI22_X1 U42 ( .A1(DATA_OUT[14]), .A2(n6), .B1(DATA_IN[14]), .B2(n2), .ZN(
        n25) );
  INV_X1 U43 ( .A(n25), .ZN(n49) );
  AOI22_X1 U44 ( .A1(DATA_OUT[15]), .A2(n6), .B1(DATA_IN[15]), .B2(n2), .ZN(
        n26) );
  INV_X1 U45 ( .A(n26), .ZN(n48) );
  AOI22_X1 U46 ( .A1(DATA_OUT[16]), .A2(n6), .B1(DATA_IN[16]), .B2(n2), .ZN(
        n27) );
  INV_X1 U47 ( .A(n27), .ZN(n47) );
  AOI22_X1 U48 ( .A1(DATA_OUT[17]), .A2(n6), .B1(DATA_IN[17]), .B2(n2), .ZN(
        n28) );
  INV_X1 U49 ( .A(n28), .ZN(n46) );
  AOI22_X1 U50 ( .A1(DATA_OUT[18]), .A2(n6), .B1(DATA_IN[18]), .B2(n2), .ZN(
        n29) );
  INV_X1 U51 ( .A(n29), .ZN(n45) );
  AOI22_X1 U52 ( .A1(DATA_OUT[19]), .A2(n6), .B1(DATA_IN[19]), .B2(n2), .ZN(
        n30) );
  INV_X1 U53 ( .A(n30), .ZN(n44) );
  AOI22_X1 U54 ( .A1(DATA_OUT[20]), .A2(n6), .B1(DATA_IN[20]), .B2(n2), .ZN(
        n31) );
  INV_X1 U55 ( .A(n31), .ZN(n43) );
  AOI22_X1 U56 ( .A1(DATA_OUT[21]), .A2(n6), .B1(DATA_IN[21]), .B2(n2), .ZN(
        n32) );
  INV_X1 U57 ( .A(n32), .ZN(n42) );
  AOI22_X1 U58 ( .A1(DATA_OUT[22]), .A2(n6), .B1(DATA_IN[22]), .B2(n2), .ZN(
        n33) );
  INV_X1 U59 ( .A(n33), .ZN(n41) );
  AOI22_X1 U60 ( .A1(DATA_OUT[23]), .A2(n6), .B1(DATA_IN[23]), .B2(n2), .ZN(
        n34) );
  INV_X1 U61 ( .A(n34), .ZN(n40) );
  AOI22_X1 U62 ( .A1(DATA_OUT[24]), .A2(n7), .B1(DATA_IN[24]), .B2(n2), .ZN(
        n35) );
  INV_X1 U63 ( .A(n35), .ZN(n39) );
  AOI22_X1 U64 ( .A1(DATA_OUT[25]), .A2(n7), .B1(DATA_IN[25]), .B2(n2), .ZN(
        n37) );
  INV_X1 U65 ( .A(n37), .ZN(n38) );
endmodule


module REG_GENERIC_NBIT5_0 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [4:0] DATA_IN;
  output [4:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n7, n8, n10, n11, n12, n13, n1, n2, n3, n4, n5, n6, n9;

  DFF_X1 \DATA_OUT_reg[4]  ( .D(n3), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n4), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n5), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n6), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n9), .CK(CLK), .Q(DATA_OUT[0]) );
  AOI22_X1 U3 ( .A1(DATA_IN[0]), .A2(n8), .B1(DATA_OUT[0]), .B2(n1), .ZN(n7)
         );
  AOI22_X1 U7 ( .A1(DATA_IN[4]), .A2(n8), .B1(DATA_OUT[4]), .B2(n1), .ZN(n13)
         );
  AOI22_X1 U6 ( .A1(DATA_IN[3]), .A2(n8), .B1(DATA_OUT[3]), .B2(n1), .ZN(n12)
         );
  AOI22_X1 U5 ( .A1(DATA_IN[2]), .A2(n8), .B1(DATA_OUT[2]), .B2(n1), .ZN(n11)
         );
  AOI22_X1 U4 ( .A1(DATA_IN[1]), .A2(n8), .B1(DATA_OUT[1]), .B2(n1), .ZN(n10)
         );
  NOR2_X1 U8 ( .A1(n2), .A2(n1), .ZN(n8) );
  NOR2_X1 U9 ( .A1(EN), .A2(n2), .ZN(n1) );
  INV_X1 U10 ( .A(RST), .ZN(n2) );
  INV_X1 U11 ( .A(n7), .ZN(n9) );
  INV_X1 U12 ( .A(n10), .ZN(n6) );
  INV_X1 U13 ( .A(n11), .ZN(n5) );
  INV_X1 U14 ( .A(n12), .ZN(n4) );
  INV_X1 U15 ( .A(n13), .ZN(n3) );
endmodule


module REG_GENERIC_NBIT5_2 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [4:0] DATA_IN;
  output [4:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  DFF_X1 \DATA_OUT_reg[4]  ( .D(n11), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n12), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n13), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n14), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n15), .CK(CLK), .Q(DATA_OUT[0]) );
  AND2_X1 U3 ( .A1(n2), .A2(n4), .ZN(n1) );
  INV_X1 U4 ( .A(n3), .ZN(n2) );
  INV_X1 U5 ( .A(RST), .ZN(n3) );
  OR2_X1 U6 ( .A1(EN), .A2(n3), .ZN(n4) );
  INV_X1 U7 ( .A(n4), .ZN(n9) );
  AOI22_X1 U8 ( .A1(DATA_OUT[0]), .A2(n9), .B1(DATA_IN[0]), .B2(n1), .ZN(n5)
         );
  INV_X1 U9 ( .A(n5), .ZN(n15) );
  AOI22_X1 U10 ( .A1(DATA_OUT[1]), .A2(n9), .B1(DATA_IN[1]), .B2(n1), .ZN(n6)
         );
  INV_X1 U11 ( .A(n6), .ZN(n14) );
  AOI22_X1 U12 ( .A1(DATA_OUT[2]), .A2(n9), .B1(DATA_IN[2]), .B2(n1), .ZN(n7)
         );
  INV_X1 U13 ( .A(n7), .ZN(n13) );
  AOI22_X1 U14 ( .A1(DATA_OUT[3]), .A2(n9), .B1(DATA_IN[3]), .B2(n1), .ZN(n8)
         );
  INV_X1 U15 ( .A(n8), .ZN(n12) );
  AOI22_X1 U16 ( .A1(DATA_OUT[4]), .A2(n9), .B1(DATA_IN[4]), .B2(n1), .ZN(n10)
         );
  INV_X1 U17 ( .A(n10), .ZN(n11) );
endmodule


module REG_GENERIC_NBIT5_1 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [4:0] DATA_IN;
  output [4:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n9, n14, n15, n16, n17, n18, n19;

  DFF_X1 \DATA_OUT_reg[4]  ( .D(n3), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n4), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n5), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n6), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n9), .CK(CLK), .Q(DATA_OUT[0]) );
  AOI22_X1 U7 ( .A1(DATA_IN[4]), .A2(n18), .B1(DATA_OUT[4]), .B2(n1), .ZN(n14)
         );
  AOI22_X1 U6 ( .A1(DATA_IN[3]), .A2(n18), .B1(DATA_OUT[3]), .B2(n1), .ZN(n15)
         );
  AOI22_X1 U5 ( .A1(DATA_IN[2]), .A2(n18), .B1(DATA_OUT[2]), .B2(n1), .ZN(n16)
         );
  AOI22_X1 U4 ( .A1(DATA_IN[1]), .A2(n18), .B1(DATA_OUT[1]), .B2(n1), .ZN(n17)
         );
  AOI22_X1 U3 ( .A1(DATA_IN[0]), .A2(n18), .B1(DATA_OUT[0]), .B2(n1), .ZN(n19)
         );
  NOR2_X1 U8 ( .A1(n2), .A2(n1), .ZN(n18) );
  NOR2_X1 U9 ( .A1(EN), .A2(n2), .ZN(n1) );
  INV_X1 U10 ( .A(RST), .ZN(n2) );
  INV_X1 U11 ( .A(n19), .ZN(n9) );
  INV_X1 U12 ( .A(n17), .ZN(n6) );
  INV_X1 U13 ( .A(n16), .ZN(n5) );
  INV_X1 U14 ( .A(n15), .ZN(n4) );
  INV_X1 U15 ( .A(n14), .ZN(n3) );
endmodule


module REG_GENERIC_NBIT32_3 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   net18836, net48248, net48246, net48244, net48254, net48252, net48250,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91;

  DFF_X1 \DATA_OUT_reg[31]  ( .D(n69), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n70), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[28]  ( .D(n19), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n71), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n72), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(net18836), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n75), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n77), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n82), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X2 \DATA_OUT_reg[13]  ( .D(n80), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X2 \DATA_OUT_reg[14]  ( .D(n79), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n78), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X2 \DATA_OUT_reg[23]  ( .D(n25), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n73), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n74), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n22), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n76), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X2 \DATA_OUT_reg[8]  ( .D(n84), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X2 \DATA_OUT_reg[7]  ( .D(n85), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X2 \DATA_OUT_reg[6]  ( .D(n86), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X2 \DATA_OUT_reg[10]  ( .D(n16), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X2 \DATA_OUT_reg[9]  ( .D(n83), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n81), .CK(CLK), .Q(DATA_OUT[12]) );
  AND2_X2 U3 ( .A1(n32), .A2(n31), .ZN(n34) );
  BUF_X1 U4 ( .A(n29), .Z(net48244) );
  OR2_X1 U5 ( .A1(n10), .A2(n35), .ZN(n13) );
  BUF_X1 U6 ( .A(n34), .Z(net48252) );
  BUF_X1 U7 ( .A(n34), .Z(net48250) );
  BUF_X1 U8 ( .A(n34), .Z(net48254) );
  NAND2_X1 U9 ( .A1(n5), .A2(n6), .ZN(n4) );
  NAND2_X1 U10 ( .A1(DATA_IN[29]), .A2(net48254), .ZN(n5) );
  OR2_X4 U11 ( .A1(n1), .A2(n10), .ZN(n6) );
  NAND2_X1 U12 ( .A1(n8), .A2(n9), .ZN(n7) );
  NAND2_X1 U13 ( .A1(net48254), .A2(DATA_IN[25]), .ZN(n8) );
  OR2_X4 U14 ( .A1(n2), .A2(n10), .ZN(n9) );
  INV_X1 U15 ( .A(n29), .ZN(n10) );
  NAND2_X1 U16 ( .A1(n12), .A2(n13), .ZN(n11) );
  NAND2_X1 U17 ( .A1(DATA_IN[0]), .A2(net48254), .ZN(n12) );
  NAND2_X1 U18 ( .A1(DATA_OUT[10]), .A2(net48244), .ZN(n14) );
  NAND2_X1 U19 ( .A1(DATA_IN[10]), .A2(net48250), .ZN(n15) );
  NAND2_X1 U20 ( .A1(n15), .A2(n14), .ZN(n16) );
  NAND2_X1 U21 ( .A1(DATA_OUT[28]), .A2(net48248), .ZN(n17) );
  NAND2_X1 U22 ( .A1(DATA_IN[28]), .A2(net48254), .ZN(n18) );
  NAND2_X1 U23 ( .A1(n18), .A2(n17), .ZN(n19) );
  NAND2_X1 U24 ( .A1(DATA_OUT[26]), .A2(net48248), .ZN(n20) );
  NAND2_X1 U25 ( .A1(DATA_IN[26]), .A2(net48254), .ZN(n21) );
  NAND2_X1 U26 ( .A1(n21), .A2(n20), .ZN(n22) );
  NAND2_X1 U27 ( .A1(DATA_OUT[23]), .A2(net48246), .ZN(n23) );
  NAND2_X1 U28 ( .A1(DATA_IN[23]), .A2(net48252), .ZN(n24) );
  NAND2_X1 U29 ( .A1(n24), .A2(n23), .ZN(n25) );
  NAND2_X1 U30 ( .A1(DATA_IN[19]), .A2(net48254), .ZN(n26) );
  OR2_X1 U31 ( .A1(n3), .A2(n10), .ZN(n27) );
  NAND2_X1 U32 ( .A1(n26), .A2(n27), .ZN(n28) );
  AOI22_X1 U33 ( .A1(DATA_IN[24]), .A2(n34), .B1(net48248), .B2(DATA_OUT[24]), 
        .ZN(n65) );
  AOI22_X1 U34 ( .A1(DATA_IN[31]), .A2(n34), .B1(net48248), .B2(DATA_OUT[31]), 
        .ZN(n68) );
  AOI22_X1 U35 ( .A1(DATA_IN[6]), .A2(n34), .B1(n29), .B2(DATA_OUT[6]), .ZN(
        n51) );
  AOI22_X1 U36 ( .A1(DATA_IN[15]), .A2(n34), .B1(net48246), .B2(DATA_OUT[15]), 
        .ZN(n59) );
  CLKBUF_X3 U37 ( .A(n29), .Z(net48246) );
  AOI22_X1 U38 ( .A1(DATA_IN[7]), .A2(n34), .B1(n29), .B2(DATA_OUT[7]), .ZN(
        n52) );
  BUF_X2 U39 ( .A(n29), .Z(net48248) );
  AOI22_X1 U40 ( .A1(DATA_IN[12]), .A2(n34), .B1(net48246), .B2(DATA_OUT[12]), 
        .ZN(n56) );
  AOI22_X1 U41 ( .A1(DATA_IN[11]), .A2(n34), .B1(n29), .B2(DATA_OUT[11]), .ZN(
        n55) );
  AOI22_X1 U42 ( .A1(DATA_IN[13]), .A2(n34), .B1(net48246), .B2(DATA_OUT[13]), 
        .ZN(n57) );
  AOI22_X1 U43 ( .A1(DATA_IN[8]), .A2(n34), .B1(n29), .B2(DATA_OUT[8]), .ZN(
        n53) );
  INV_X2 U44 ( .A(n31), .ZN(n29) );
  AOI22_X1 U45 ( .A1(DATA_IN[9]), .A2(n34), .B1(net48244), .B2(DATA_OUT[9]), 
        .ZN(n54) );
  AOI22_X1 U46 ( .A1(DATA_IN[27]), .A2(n34), .B1(net48248), .B2(DATA_OUT[27]), 
        .ZN(n66) );
  AOI22_X1 U47 ( .A1(DATA_IN[30]), .A2(n34), .B1(net48248), .B2(DATA_OUT[30]), 
        .ZN(n67) );
  AOI22_X1 U48 ( .A1(DATA_IN[22]), .A2(n34), .B1(net48246), .B2(DATA_OUT[22]), 
        .ZN(n30) );
  INV_X1 U49 ( .A(n30), .ZN(net18836) );
  INV_X1 U50 ( .A(n33), .ZN(n32) );
  INV_X1 U51 ( .A(RST), .ZN(n33) );
  OR2_X1 U52 ( .A1(n33), .A2(EN), .ZN(n31) );
  AOI22_X1 U58 ( .A1(DATA_OUT[1]), .A2(net48244), .B1(DATA_IN[1]), .B2(
        net48250), .ZN(n46) );
  INV_X1 U59 ( .A(n46), .ZN(n91) );
  AOI22_X1 U60 ( .A1(DATA_OUT[2]), .A2(net48244), .B1(DATA_IN[2]), .B2(
        net48250), .ZN(n47) );
  INV_X1 U61 ( .A(n47), .ZN(n90) );
  AOI22_X1 U62 ( .A1(DATA_OUT[3]), .A2(net48244), .B1(DATA_IN[3]), .B2(
        net48250), .ZN(n48) );
  INV_X1 U63 ( .A(n48), .ZN(n89) );
  AOI22_X1 U64 ( .A1(DATA_OUT[4]), .A2(net48244), .B1(DATA_IN[4]), .B2(
        net48250), .ZN(n49) );
  INV_X1 U65 ( .A(n49), .ZN(n88) );
  AOI22_X1 U66 ( .A1(DATA_OUT[5]), .A2(net48244), .B1(DATA_IN[5]), .B2(
        net48250), .ZN(n50) );
  INV_X1 U67 ( .A(n50), .ZN(n87) );
  INV_X1 U68 ( .A(n51), .ZN(n86) );
  INV_X1 U69 ( .A(n52), .ZN(n85) );
  INV_X1 U70 ( .A(n53), .ZN(n84) );
  INV_X1 U71 ( .A(n54), .ZN(n83) );
  INV_X1 U72 ( .A(n55), .ZN(n82) );
  INV_X1 U73 ( .A(n56), .ZN(n81) );
  INV_X1 U74 ( .A(n57), .ZN(n80) );
  AOI22_X1 U75 ( .A1(DATA_OUT[14]), .A2(net48246), .B1(DATA_IN[14]), .B2(
        net48252), .ZN(n58) );
  INV_X1 U76 ( .A(n58), .ZN(n79) );
  INV_X1 U77 ( .A(n59), .ZN(n78) );
  AOI22_X1 U78 ( .A1(DATA_OUT[16]), .A2(net48246), .B1(DATA_IN[16]), .B2(
        net48252), .ZN(n60) );
  INV_X1 U79 ( .A(n60), .ZN(n77) );
  AOI22_X1 U80 ( .A1(DATA_OUT[17]), .A2(net48246), .B1(DATA_IN[17]), .B2(
        net48252), .ZN(n61) );
  INV_X1 U81 ( .A(n61), .ZN(n76) );
  AOI22_X1 U82 ( .A1(DATA_OUT[18]), .A2(net48246), .B1(DATA_IN[18]), .B2(
        net48252), .ZN(n62) );
  INV_X1 U83 ( .A(n62), .ZN(n75) );
  AOI22_X1 U84 ( .A1(DATA_OUT[20]), .A2(net48246), .B1(DATA_IN[20]), .B2(
        net48252), .ZN(n63) );
  INV_X1 U85 ( .A(n63), .ZN(n74) );
  AOI22_X1 U86 ( .A1(DATA_OUT[21]), .A2(net48246), .B1(DATA_IN[21]), .B2(
        net48252), .ZN(n64) );
  INV_X1 U87 ( .A(n64), .ZN(n73) );
  INV_X1 U88 ( .A(n65), .ZN(n72) );
  INV_X1 U89 ( .A(n66), .ZN(n71) );
  INV_X1 U90 ( .A(n67), .ZN(n70) );
  INV_X1 U91 ( .A(n68), .ZN(n69) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n11), .CK(CLK), .Q(DATA_OUT[0]), .QN(n35) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n4), .CK(CLK), .Q(DATA_OUT[29]), .QN(n1) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n91), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n90), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n87), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n88), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n89), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n28), .CK(CLK), .Q(DATA_OUT[19]), .QN(n3) );
  DFF_X1 \DATA_OUT_reg[25]  ( .D(n7), .CK(CLK), .Q(DATA_OUT[25]), .QN(n2) );
endmodule


module REG_GENERIC_NBIT32_2 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139;

  BUF_X2 U35 ( .A(n106), .Z(n69) );
  BUF_X2 U36 ( .A(n106), .Z(n70) );
  BUF_X1 U37 ( .A(n65), .Z(n66) );
  BUF_X1 U38 ( .A(n65), .Z(n67) );
  BUF_X2 U39 ( .A(n106), .Z(n71) );
  BUF_X1 U40 ( .A(n65), .Z(n68) );
  AND2_X1 U41 ( .A1(n72), .A2(n74), .ZN(n65) );
  INV_X1 U42 ( .A(n73), .ZN(n72) );
  INV_X1 U43 ( .A(RST), .ZN(n73) );
  OR2_X1 U44 ( .A1(EN), .A2(n73), .ZN(n74) );
  INV_X1 U45 ( .A(n74), .ZN(n106) );
  AOI22_X1 U46 ( .A1(DATA_OUT[0]), .A2(n69), .B1(DATA_IN[0]), .B2(n66), .ZN(
        n75) );
  INV_X1 U47 ( .A(n75), .ZN(n139) );
  AOI22_X1 U48 ( .A1(DATA_OUT[1]), .A2(n69), .B1(DATA_IN[1]), .B2(n66), .ZN(
        n76) );
  INV_X1 U49 ( .A(n76), .ZN(n138) );
  AOI22_X1 U50 ( .A1(DATA_OUT[2]), .A2(n69), .B1(DATA_IN[2]), .B2(n66), .ZN(
        n77) );
  INV_X1 U51 ( .A(n77), .ZN(n137) );
  AOI22_X1 U52 ( .A1(DATA_OUT[3]), .A2(n69), .B1(DATA_IN[3]), .B2(n66), .ZN(
        n78) );
  INV_X1 U53 ( .A(n78), .ZN(n136) );
  AOI22_X1 U54 ( .A1(DATA_OUT[4]), .A2(n69), .B1(DATA_IN[4]), .B2(n66), .ZN(
        n79) );
  INV_X1 U55 ( .A(n79), .ZN(n135) );
  AOI22_X1 U56 ( .A1(DATA_OUT[5]), .A2(n69), .B1(DATA_IN[5]), .B2(n66), .ZN(
        n80) );
  INV_X1 U57 ( .A(n80), .ZN(n134) );
  AOI22_X1 U58 ( .A1(DATA_OUT[6]), .A2(n69), .B1(DATA_IN[6]), .B2(n66), .ZN(
        n81) );
  INV_X1 U59 ( .A(n81), .ZN(n133) );
  AOI22_X1 U60 ( .A1(DATA_OUT[7]), .A2(n69), .B1(DATA_IN[7]), .B2(n66), .ZN(
        n82) );
  INV_X1 U61 ( .A(n82), .ZN(n132) );
  AOI22_X1 U62 ( .A1(DATA_OUT[8]), .A2(n69), .B1(DATA_IN[8]), .B2(n66), .ZN(
        n83) );
  INV_X1 U63 ( .A(n83), .ZN(n131) );
  AOI22_X1 U64 ( .A1(DATA_OUT[9]), .A2(n69), .B1(DATA_IN[9]), .B2(n66), .ZN(
        n84) );
  INV_X1 U65 ( .A(n84), .ZN(n130) );
  AOI22_X1 U66 ( .A1(DATA_OUT[10]), .A2(n69), .B1(DATA_IN[10]), .B2(n66), .ZN(
        n85) );
  INV_X1 U67 ( .A(n85), .ZN(n129) );
  AOI22_X1 U68 ( .A1(DATA_OUT[11]), .A2(n69), .B1(DATA_IN[11]), .B2(n66), .ZN(
        n86) );
  INV_X1 U69 ( .A(n86), .ZN(n128) );
  AOI22_X1 U70 ( .A1(DATA_OUT[12]), .A2(n70), .B1(DATA_IN[12]), .B2(n67), .ZN(
        n87) );
  INV_X1 U71 ( .A(n87), .ZN(n127) );
  AOI22_X1 U72 ( .A1(DATA_OUT[13]), .A2(n70), .B1(DATA_IN[13]), .B2(n67), .ZN(
        n88) );
  INV_X1 U73 ( .A(n88), .ZN(n126) );
  AOI22_X1 U74 ( .A1(DATA_OUT[14]), .A2(n70), .B1(DATA_IN[14]), .B2(n67), .ZN(
        n89) );
  INV_X1 U75 ( .A(n89), .ZN(n125) );
  AOI22_X1 U76 ( .A1(DATA_OUT[15]), .A2(n70), .B1(DATA_IN[15]), .B2(n67), .ZN(
        n90) );
  INV_X1 U77 ( .A(n90), .ZN(n124) );
  AOI22_X1 U78 ( .A1(DATA_OUT[16]), .A2(n70), .B1(DATA_IN[16]), .B2(n67), .ZN(
        n91) );
  INV_X1 U79 ( .A(n91), .ZN(n123) );
  AOI22_X1 U80 ( .A1(DATA_OUT[17]), .A2(n70), .B1(DATA_IN[17]), .B2(n67), .ZN(
        n92) );
  INV_X1 U81 ( .A(n92), .ZN(n122) );
  AOI22_X1 U82 ( .A1(DATA_OUT[18]), .A2(n70), .B1(DATA_IN[18]), .B2(n67), .ZN(
        n93) );
  INV_X1 U83 ( .A(n93), .ZN(n121) );
  AOI22_X1 U84 ( .A1(DATA_OUT[19]), .A2(n70), .B1(DATA_IN[19]), .B2(n67), .ZN(
        n94) );
  INV_X1 U85 ( .A(n94), .ZN(n120) );
  AOI22_X1 U86 ( .A1(DATA_OUT[20]), .A2(n70), .B1(DATA_IN[20]), .B2(n67), .ZN(
        n95) );
  INV_X1 U87 ( .A(n95), .ZN(n119) );
  AOI22_X1 U88 ( .A1(DATA_OUT[21]), .A2(n70), .B1(DATA_IN[21]), .B2(n67), .ZN(
        n96) );
  INV_X1 U89 ( .A(n96), .ZN(n118) );
  AOI22_X1 U90 ( .A1(DATA_OUT[22]), .A2(n70), .B1(DATA_IN[22]), .B2(n67), .ZN(
        n97) );
  INV_X1 U91 ( .A(n97), .ZN(n117) );
  AOI22_X1 U92 ( .A1(DATA_OUT[23]), .A2(n70), .B1(DATA_IN[23]), .B2(n67), .ZN(
        n98) );
  INV_X1 U93 ( .A(n98), .ZN(n116) );
  AOI22_X1 U94 ( .A1(DATA_OUT[24]), .A2(n71), .B1(DATA_IN[24]), .B2(n68), .ZN(
        n99) );
  INV_X1 U95 ( .A(n99), .ZN(n115) );
  AOI22_X1 U96 ( .A1(DATA_OUT[25]), .A2(n71), .B1(DATA_IN[25]), .B2(n68), .ZN(
        n100) );
  INV_X1 U97 ( .A(n100), .ZN(n114) );
  AOI22_X1 U98 ( .A1(DATA_OUT[26]), .A2(n71), .B1(DATA_IN[26]), .B2(n68), .ZN(
        n101) );
  INV_X1 U99 ( .A(n101), .ZN(n113) );
  AOI22_X1 U100 ( .A1(DATA_OUT[27]), .A2(n71), .B1(DATA_IN[27]), .B2(n68), 
        .ZN(n102) );
  INV_X1 U101 ( .A(n102), .ZN(n112) );
  AOI22_X1 U102 ( .A1(DATA_OUT[28]), .A2(n71), .B1(DATA_IN[28]), .B2(n68), 
        .ZN(n103) );
  INV_X1 U103 ( .A(n103), .ZN(n111) );
  AOI22_X1 U104 ( .A1(DATA_OUT[29]), .A2(n71), .B1(DATA_IN[29]), .B2(n68), 
        .ZN(n104) );
  INV_X1 U105 ( .A(n104), .ZN(n110) );
  AOI22_X1 U106 ( .A1(DATA_OUT[30]), .A2(n71), .B1(DATA_IN[30]), .B2(n68), 
        .ZN(n105) );
  INV_X1 U107 ( .A(n105), .ZN(n109) );
  AOI22_X1 U108 ( .A1(DATA_OUT[31]), .A2(n71), .B1(DATA_IN[31]), .B2(n68), 
        .ZN(n107) );
  INV_X1 U109 ( .A(n107), .ZN(n108) );
  DFF_X1 \DATA_OUT_reg[31]  ( .D(n108), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n109), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n110), .CK(CLK), .Q(DATA_OUT[29]) );
  DFF_X1 \DATA_OUT_reg[28]  ( .D(n111), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n112), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n113), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[25]  ( .D(n114), .CK(CLK), .Q(DATA_OUT[25]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n115), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[23]  ( .D(n116), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n117), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n118), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n119), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n120), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n121), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n122), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n123), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n124), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n125), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n126), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n127), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n128), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n129), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n130), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n131), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n132), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n133), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n134), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n135), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n136), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n137), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n138), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n139), .CK(CLK), .Q(DATA_OUT[0]) );
endmodule


module REG_GENERIC_NBIT32_1 ( CLK, RST, EN, DATA_IN, DATA_OUT );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input CLK, RST, EN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n36, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106;

  DFF_X1 \DATA_OUT_reg[31]  ( .D(n9), .CK(CLK), .Q(DATA_OUT[31]) );
  DFF_X1 \DATA_OUT_reg[30]  ( .D(n10), .CK(CLK), .Q(DATA_OUT[30]) );
  DFF_X1 \DATA_OUT_reg[29]  ( .D(n11), .CK(CLK), .Q(DATA_OUT[29]) );
  DFF_X1 \DATA_OUT_reg[28]  ( .D(n12), .CK(CLK), .Q(DATA_OUT[28]) );
  DFF_X1 \DATA_OUT_reg[27]  ( .D(n13), .CK(CLK), .Q(DATA_OUT[27]) );
  DFF_X1 \DATA_OUT_reg[26]  ( .D(n14), .CK(CLK), .Q(DATA_OUT[26]) );
  DFF_X1 \DATA_OUT_reg[25]  ( .D(n15), .CK(CLK), .Q(DATA_OUT[25]) );
  DFF_X1 \DATA_OUT_reg[24]  ( .D(n16), .CK(CLK), .Q(DATA_OUT[24]) );
  DFF_X1 \DATA_OUT_reg[23]  ( .D(n17), .CK(CLK), .Q(DATA_OUT[23]) );
  DFF_X1 \DATA_OUT_reg[22]  ( .D(n18), .CK(CLK), .Q(DATA_OUT[22]) );
  DFF_X1 \DATA_OUT_reg[21]  ( .D(n19), .CK(CLK), .Q(DATA_OUT[21]) );
  DFF_X1 \DATA_OUT_reg[20]  ( .D(n20), .CK(CLK), .Q(DATA_OUT[20]) );
  DFF_X1 \DATA_OUT_reg[19]  ( .D(n21), .CK(CLK), .Q(DATA_OUT[19]) );
  DFF_X1 \DATA_OUT_reg[18]  ( .D(n22), .CK(CLK), .Q(DATA_OUT[18]) );
  DFF_X1 \DATA_OUT_reg[17]  ( .D(n23), .CK(CLK), .Q(DATA_OUT[17]) );
  DFF_X1 \DATA_OUT_reg[16]  ( .D(n24), .CK(CLK), .Q(DATA_OUT[16]) );
  DFF_X1 \DATA_OUT_reg[15]  ( .D(n25), .CK(CLK), .Q(DATA_OUT[15]) );
  DFF_X1 \DATA_OUT_reg[14]  ( .D(n26), .CK(CLK), .Q(DATA_OUT[14]) );
  DFF_X1 \DATA_OUT_reg[13]  ( .D(n27), .CK(CLK), .Q(DATA_OUT[13]) );
  DFF_X1 \DATA_OUT_reg[12]  ( .D(n28), .CK(CLK), .Q(DATA_OUT[12]) );
  DFF_X1 \DATA_OUT_reg[11]  ( .D(n29), .CK(CLK), .Q(DATA_OUT[11]) );
  DFF_X1 \DATA_OUT_reg[10]  ( .D(n30), .CK(CLK), .Q(DATA_OUT[10]) );
  DFF_X1 \DATA_OUT_reg[9]  ( .D(n31), .CK(CLK), .Q(DATA_OUT[9]) );
  DFF_X1 \DATA_OUT_reg[8]  ( .D(n32), .CK(CLK), .Q(DATA_OUT[8]) );
  DFF_X1 \DATA_OUT_reg[7]  ( .D(n33), .CK(CLK), .Q(DATA_OUT[7]) );
  DFF_X1 \DATA_OUT_reg[6]  ( .D(n36), .CK(CLK), .Q(DATA_OUT[6]) );
  DFF_X1 \DATA_OUT_reg[5]  ( .D(n68), .CK(CLK), .Q(DATA_OUT[5]) );
  DFF_X1 \DATA_OUT_reg[4]  ( .D(n69), .CK(CLK), .Q(DATA_OUT[4]) );
  DFF_X1 \DATA_OUT_reg[3]  ( .D(n70), .CK(CLK), .Q(DATA_OUT[3]) );
  DFF_X1 \DATA_OUT_reg[2]  ( .D(n71), .CK(CLK), .Q(DATA_OUT[2]) );
  DFF_X1 \DATA_OUT_reg[1]  ( .D(n72), .CK(CLK), .Q(DATA_OUT[1]) );
  DFF_X1 \DATA_OUT_reg[0]  ( .D(n73), .CK(CLK), .Q(DATA_OUT[0]) );
  AOI22_X1 U25 ( .A1(DATA_IN[22]), .A2(n5), .B1(DATA_OUT[22]), .B2(n3), .ZN(
        n83) );
  AOI22_X1 U9 ( .A1(DATA_IN[6]), .A2(n7), .B1(DATA_OUT[6]), .B2(n2), .ZN(n99)
         );
  AOI22_X1 U8 ( .A1(DATA_IN[5]), .A2(n7), .B1(DATA_OUT[5]), .B2(n2), .ZN(n100)
         );
  AOI22_X1 U7 ( .A1(DATA_IN[4]), .A2(n7), .B1(DATA_OUT[4]), .B2(n2), .ZN(n101)
         );
  AOI22_X1 U6 ( .A1(DATA_IN[3]), .A2(n7), .B1(DATA_OUT[3]), .B2(n2), .ZN(n102)
         );
  AOI22_X1 U5 ( .A1(DATA_IN[2]), .A2(n7), .B1(DATA_OUT[2]), .B2(n2), .ZN(n103)
         );
  AOI22_X1 U4 ( .A1(DATA_IN[1]), .A2(n7), .B1(DATA_OUT[1]), .B2(n2), .ZN(n104)
         );
  AOI22_X1 U3 ( .A1(DATA_IN[0]), .A2(n7), .B1(DATA_OUT[0]), .B2(n2), .ZN(n106)
         );
  AOI22_X1 U10 ( .A1(DATA_IN[7]), .A2(n7), .B1(DATA_OUT[7]), .B2(n2), .ZN(n98)
         );
  AOI22_X1 U34 ( .A1(DATA_IN[31]), .A2(n5), .B1(DATA_OUT[31]), .B2(n4), .ZN(
        n74) );
  AOI22_X1 U33 ( .A1(DATA_IN[30]), .A2(n5), .B1(DATA_OUT[30]), .B2(n4), .ZN(
        n75) );
  AOI22_X1 U32 ( .A1(DATA_IN[29]), .A2(n5), .B1(DATA_OUT[29]), .B2(n4), .ZN(
        n76) );
  AOI22_X1 U31 ( .A1(DATA_IN[28]), .A2(n5), .B1(DATA_OUT[28]), .B2(n4), .ZN(
        n77) );
  AOI22_X1 U30 ( .A1(DATA_IN[27]), .A2(n5), .B1(DATA_OUT[27]), .B2(n4), .ZN(
        n78) );
  AOI22_X1 U29 ( .A1(DATA_IN[26]), .A2(n5), .B1(DATA_OUT[26]), .B2(n4), .ZN(
        n79) );
  AOI22_X1 U28 ( .A1(DATA_IN[25]), .A2(n5), .B1(DATA_OUT[25]), .B2(n4), .ZN(
        n80) );
  AOI22_X1 U27 ( .A1(DATA_IN[24]), .A2(n5), .B1(DATA_OUT[24]), .B2(n4), .ZN(
        n81) );
  AOI22_X1 U26 ( .A1(DATA_IN[23]), .A2(n5), .B1(DATA_OUT[23]), .B2(n3), .ZN(
        n82) );
  AOI22_X1 U24 ( .A1(DATA_IN[21]), .A2(n5), .B1(DATA_OUT[21]), .B2(n3), .ZN(
        n84) );
  AOI22_X1 U23 ( .A1(DATA_IN[20]), .A2(n5), .B1(DATA_OUT[20]), .B2(n3), .ZN(
        n85) );
  AOI22_X1 U22 ( .A1(DATA_IN[19]), .A2(n6), .B1(DATA_OUT[19]), .B2(n3), .ZN(
        n86) );
  AOI22_X1 U21 ( .A1(DATA_IN[18]), .A2(n6), .B1(DATA_OUT[18]), .B2(n3), .ZN(
        n87) );
  AOI22_X1 U20 ( .A1(DATA_IN[17]), .A2(n6), .B1(DATA_OUT[17]), .B2(n3), .ZN(
        n88) );
  AOI22_X1 U19 ( .A1(DATA_IN[16]), .A2(n6), .B1(DATA_OUT[16]), .B2(n3), .ZN(
        n89) );
  AOI22_X1 U18 ( .A1(DATA_IN[15]), .A2(n6), .B1(DATA_OUT[15]), .B2(n3), .ZN(
        n90) );
  AOI22_X1 U17 ( .A1(DATA_IN[14]), .A2(n6), .B1(DATA_OUT[14]), .B2(n3), .ZN(
        n91) );
  AOI22_X1 U16 ( .A1(DATA_IN[13]), .A2(n6), .B1(DATA_OUT[13]), .B2(n3), .ZN(
        n92) );
  AOI22_X1 U15 ( .A1(DATA_IN[12]), .A2(n6), .B1(DATA_OUT[12]), .B2(n3), .ZN(
        n93) );
  AOI22_X1 U14 ( .A1(DATA_IN[11]), .A2(n6), .B1(DATA_OUT[11]), .B2(n2), .ZN(
        n94) );
  AOI22_X1 U13 ( .A1(DATA_IN[10]), .A2(n6), .B1(DATA_OUT[10]), .B2(n2), .ZN(
        n95) );
  AOI22_X1 U12 ( .A1(DATA_IN[9]), .A2(n6), .B1(DATA_OUT[9]), .B2(n2), .ZN(n96)
         );
  AOI22_X1 U11 ( .A1(DATA_IN[8]), .A2(n6), .B1(DATA_OUT[8]), .B2(n2), .ZN(n97)
         );
  NOR2_X1 U35 ( .A1(n8), .A2(n4), .ZN(n105) );
  BUF_X2 U36 ( .A(n105), .Z(n6) );
  BUF_X1 U37 ( .A(n105), .Z(n7) );
  BUF_X2 U38 ( .A(n105), .Z(n5) );
  BUF_X1 U39 ( .A(n1), .Z(n3) );
  BUF_X1 U40 ( .A(n1), .Z(n2) );
  BUF_X1 U41 ( .A(n1), .Z(n4) );
  NOR2_X1 U42 ( .A1(EN), .A2(n8), .ZN(n1) );
  INV_X1 U43 ( .A(RST), .ZN(n8) );
  INV_X1 U44 ( .A(n106), .ZN(n73) );
  INV_X1 U45 ( .A(n104), .ZN(n72) );
  INV_X1 U46 ( .A(n103), .ZN(n71) );
  INV_X1 U47 ( .A(n102), .ZN(n70) );
  INV_X1 U48 ( .A(n101), .ZN(n69) );
  INV_X1 U49 ( .A(n100), .ZN(n68) );
  INV_X1 U50 ( .A(n99), .ZN(n36) );
  INV_X1 U51 ( .A(n98), .ZN(n33) );
  INV_X1 U52 ( .A(n97), .ZN(n32) );
  INV_X1 U53 ( .A(n96), .ZN(n31) );
  INV_X1 U54 ( .A(n95), .ZN(n30) );
  INV_X1 U55 ( .A(n94), .ZN(n29) );
  INV_X1 U56 ( .A(n93), .ZN(n28) );
  INV_X1 U57 ( .A(n92), .ZN(n27) );
  INV_X1 U58 ( .A(n91), .ZN(n26) );
  INV_X1 U59 ( .A(n90), .ZN(n25) );
  INV_X1 U60 ( .A(n89), .ZN(n24) );
  INV_X1 U61 ( .A(n88), .ZN(n23) );
  INV_X1 U62 ( .A(n87), .ZN(n22) );
  INV_X1 U63 ( .A(n86), .ZN(n21) );
  INV_X1 U64 ( .A(n85), .ZN(n20) );
  INV_X1 U65 ( .A(n84), .ZN(n19) );
  INV_X1 U66 ( .A(n83), .ZN(n18) );
  INV_X1 U67 ( .A(n82), .ZN(n17) );
  INV_X1 U68 ( .A(n81), .ZN(n16) );
  INV_X1 U69 ( .A(n80), .ZN(n15) );
  INV_X1 U70 ( .A(n79), .ZN(n14) );
  INV_X1 U71 ( .A(n78), .ZN(n13) );
  INV_X1 U72 ( .A(n77), .ZN(n12) );
  INV_X1 U73 ( .A(n76), .ZN(n11) );
  INV_X1 U74 ( .A(n75), .ZN(n10) );
  INV_X1 U75 ( .A(n74), .ZN(n9) );
endmodule


module BRANCHING_UNIT_N32 ( CLK, RST, Reg_A, EQ_cond, IS_JUMP, branch_taken );
  input [31:0] Reg_A;
  input CLK, RST, EQ_cond, IS_JUMP;
  output branch_taken;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  DFF_X1 branch_taken_reg ( .D(n14), .CK(CLK), .Q(branch_taken) );
  NOR4_X1 U3 ( .A1(Reg_A[19]), .A2(Reg_A[18]), .A3(Reg_A[17]), .A4(Reg_A[16]), 
        .ZN(n4) );
  NOR4_X1 U4 ( .A1(Reg_A[23]), .A2(Reg_A[22]), .A3(Reg_A[21]), .A4(Reg_A[20]), 
        .ZN(n3) );
  NOR4_X1 U5 ( .A1(Reg_A[27]), .A2(Reg_A[26]), .A3(Reg_A[25]), .A4(Reg_A[24]), 
        .ZN(n2) );
  NOR4_X1 U6 ( .A1(Reg_A[31]), .A2(Reg_A[30]), .A3(Reg_A[29]), .A4(Reg_A[28]), 
        .ZN(n1) );
  NAND4_X1 U7 ( .A1(n4), .A2(n3), .A3(n2), .A4(n1), .ZN(n10) );
  NOR4_X1 U8 ( .A1(Reg_A[3]), .A2(Reg_A[2]), .A3(Reg_A[1]), .A4(Reg_A[0]), 
        .ZN(n8) );
  NOR4_X1 U9 ( .A1(Reg_A[7]), .A2(Reg_A[6]), .A3(Reg_A[5]), .A4(Reg_A[4]), 
        .ZN(n7) );
  NOR4_X1 U10 ( .A1(Reg_A[11]), .A2(Reg_A[10]), .A3(Reg_A[9]), .A4(Reg_A[8]), 
        .ZN(n6) );
  NOR4_X1 U11 ( .A1(Reg_A[15]), .A2(Reg_A[14]), .A3(Reg_A[13]), .A4(Reg_A[12]), 
        .ZN(n5) );
  NAND4_X1 U12 ( .A1(n8), .A2(n7), .A3(n6), .A4(n5), .ZN(n9) );
  NOR2_X1 U13 ( .A1(n10), .A2(n9), .ZN(n11) );
  XNOR2_X1 U14 ( .A(EQ_cond), .B(n11), .ZN(n12) );
  OAI21_X1 U15 ( .B1(IS_JUMP), .B2(n12), .A(RST), .ZN(n13) );
  INV_X1 U16 ( .A(n13), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  BUF_X2 U1 ( .A(SEL), .Z(n1) );
  BUF_X2 U2 ( .A(SEL), .Z(n3) );
  BUF_X2 U3 ( .A(SEL), .Z(n2) );
  MUX2_X1 U4 ( .A(A[0]), .B(B[0]), .S(n3), .Z(Y[0]) );
  MUX2_X1 U5 ( .A(A[1]), .B(B[1]), .S(n2), .Z(Y[1]) );
  MUX2_X1 U6 ( .A(A[2]), .B(B[2]), .S(n2), .Z(Y[2]) );
  MUX2_X1 U7 ( .A(A[3]), .B(B[3]), .S(n2), .Z(Y[3]) );
  MUX2_X1 U8 ( .A(A[4]), .B(B[4]), .S(n2), .Z(Y[4]) );
  MUX2_X1 U9 ( .A(A[5]), .B(B[5]), .S(n3), .Z(Y[5]) );
  MUX2_X1 U10 ( .A(A[6]), .B(B[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U11 ( .A(A[7]), .B(B[7]), .S(n3), .Z(Y[7]) );
  MUX2_X1 U12 ( .A(A[8]), .B(B[8]), .S(n1), .Z(Y[8]) );
  MUX2_X1 U13 ( .A(A[9]), .B(B[9]), .S(n1), .Z(Y[9]) );
  MUX2_X1 U14 ( .A(A[10]), .B(B[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U15 ( .A(A[11]), .B(B[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U16 ( .A(A[12]), .B(B[12]), .S(n3), .Z(Y[12]) );
  MUX2_X1 U17 ( .A(A[13]), .B(B[13]), .S(n1), .Z(Y[13]) );
  MUX2_X1 U18 ( .A(A[14]), .B(B[14]), .S(n3), .Z(Y[14]) );
  MUX2_X1 U19 ( .A(A[15]), .B(B[15]), .S(n3), .Z(Y[15]) );
  MUX2_X1 U20 ( .A(A[16]), .B(B[16]), .S(n2), .Z(Y[16]) );
  MUX2_X1 U21 ( .A(A[17]), .B(B[17]), .S(n3), .Z(Y[17]) );
  MUX2_X1 U22 ( .A(A[18]), .B(B[18]), .S(n2), .Z(Y[18]) );
  MUX2_X1 U23 ( .A(A[19]), .B(B[19]), .S(n2), .Z(Y[19]) );
  MUX2_X1 U24 ( .A(A[20]), .B(B[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U25 ( .A(A[21]), .B(B[21]), .S(n3), .Z(Y[21]) );
  MUX2_X1 U26 ( .A(A[22]), .B(B[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U27 ( .A(A[23]), .B(B[23]), .S(n3), .Z(Y[23]) );
  MUX2_X1 U28 ( .A(A[24]), .B(B[24]), .S(n3), .Z(Y[24]) );
  MUX2_X1 U29 ( .A(A[25]), .B(B[25]), .S(n3), .Z(Y[25]) );
  MUX2_X1 U30 ( .A(A[26]), .B(B[26]), .S(n2), .Z(Y[26]) );
  MUX2_X1 U31 ( .A(A[27]), .B(B[27]), .S(n2), .Z(Y[27]) );
  MUX2_X1 U32 ( .A(A[28]), .B(B[28]), .S(n3), .Z(Y[28]) );
  MUX2_X1 U33 ( .A(A[29]), .B(B[29]), .S(n2), .Z(Y[29]) );
  MUX2_X1 U34 ( .A(A[30]), .B(B[30]), .S(n3), .Z(Y[30]) );
  MUX2_X1 U35 ( .A(A[31]), .B(B[31]), .S(n2), .Z(Y[31]) );
endmodule


module MUX21 ( A, B, SEL, Y );
  input A, B, SEL;
  output Y;


  MUX2_X1 U1 ( .A(A), .B(B), .S(SEL), .Z(Y) );
endmodule


module MUX21_GENERIC_NBIT5_0 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(A[0]), .B(B[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(A[1]), .B(B[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(A[2]), .B(B[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(A[3]), .B(B[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U5 ( .A(A[4]), .B(B[4]), .S(SEL), .Z(Y[4]) );
endmodule


module MUX21_GENERIC_NBIT32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   net19168, net47414, net47410, net47408, net52261, net52463, net52635,
         net52857, net52936, net52945, n1, n2, n3, n4, n5, n6, n8, n9, n10,
         n11, n12, n14, n15, n16, n17, n18, n19, n20, n21;
  assign Y[12] = net19168;

  MUX2_X2 U1 ( .A(B[30]), .B(A[30]), .S(n9), .Z(Y[30]) );
  INV_X1 U2 ( .A(n14), .ZN(n1) );
  INV_X1 U3 ( .A(n14), .ZN(net52945) );
  OR2_X2 U4 ( .A1(n5), .A2(n6), .ZN(Y[21]) );
  MUX2_X1 U5 ( .A(A[24]), .B(B[24]), .S(n3), .Z(Y[24]) );
  MUX2_X1 U6 ( .A(A[29]), .B(B[29]), .S(n3), .Z(Y[29]) );
  CLKBUF_X1 U7 ( .A(net47414), .Z(n2) );
  INV_X1 U8 ( .A(net47414), .ZN(net52463) );
  INV_X1 U9 ( .A(net47414), .ZN(n3) );
  INV_X1 U10 ( .A(A[21]), .ZN(n4) );
  NOR2_X1 U11 ( .A1(n3), .A2(n4), .ZN(n6) );
  AND2_X1 U12 ( .A1(B[21]), .A2(net52261), .ZN(n5) );
  INV_X1 U13 ( .A(B[18]), .ZN(n8) );
  INV_X1 U14 ( .A(net52945), .ZN(n9) );
  INV_X1 U15 ( .A(A[18]), .ZN(n10) );
  NOR2_X1 U16 ( .A1(n8), .A2(n9), .ZN(n11) );
  NOR2_X1 U17 ( .A1(net52463), .A2(n10), .ZN(n12) );
  OR2_X4 U18 ( .A1(n11), .A2(n12), .ZN(Y[18]) );
  MUX2_X1 U19 ( .A(B[5]), .B(A[5]), .S(net52936), .Z(Y[5]) );
  MUX2_X1 U20 ( .A(A[12]), .B(B[12]), .S(net47408), .Z(net19168) );
  INV_X1 U21 ( .A(SEL), .ZN(n14) );
  INV_X1 U22 ( .A(n14), .ZN(net52261) );
  INV_X1 U23 ( .A(n14), .ZN(net47410) );
  BUF_X1 U24 ( .A(SEL), .Z(net52635) );
  INV_X1 U25 ( .A(SEL), .ZN(net47414) );
  MUX2_X1 U26 ( .A(A[19]), .B(B[19]), .S(net52463), .Z(Y[19]) );
  INV_X1 U27 ( .A(net47410), .ZN(net52936) );
  MUX2_X1 U28 ( .A(A[16]), .B(B[16]), .S(net52945), .Z(Y[16]) );
  NAND2_X1 U29 ( .A1(A[15]), .A2(net52857), .ZN(n15) );
  NAND2_X1 U30 ( .A1(B[15]), .A2(net52261), .ZN(n16) );
  NAND2_X2 U31 ( .A1(n15), .A2(n16), .ZN(Y[15]) );
  INV_X1 U32 ( .A(n1), .ZN(net52857) );
  INV_X2 U33 ( .A(n21), .ZN(Y[2]) );
  INV_X1 U34 ( .A(net47414), .ZN(net47408) );
  MUX2_X1 U35 ( .A(B[13]), .B(A[13]), .S(net47414), .Z(Y[13]) );
  NAND2_X1 U36 ( .A1(n17), .A2(n18), .ZN(Y[3]) );
  MUX2_X1 U37 ( .A(A[14]), .B(B[14]), .S(n1), .Z(Y[14]) );
  NAND2_X1 U38 ( .A1(A[3]), .A2(n2), .ZN(n17) );
  NAND2_X1 U39 ( .A1(B[3]), .A2(net52945), .ZN(n18) );
  MUX2_X1 U40 ( .A(A[7]), .B(B[7]), .S(net47410), .Z(Y[7]) );
  MUX2_X1 U41 ( .A(A[8]), .B(B[8]), .S(net52635), .Z(Y[8]) );
  AOI22_X1 U42 ( .A1(A[0]), .A2(n2), .B1(B[0]), .B2(net52945), .ZN(n19) );
  INV_X1 U43 ( .A(n19), .ZN(Y[0]) );
  AOI22_X1 U44 ( .A1(net52261), .A2(B[1]), .B1(net47414), .B2(A[1]), .ZN(n20)
         );
  INV_X1 U45 ( .A(n20), .ZN(Y[1]) );
  AOI22_X1 U46 ( .A1(net47414), .A2(A[2]), .B1(net52635), .B2(B[2]), .ZN(n21)
         );
  MUX2_X1 U47 ( .A(A[4]), .B(B[4]), .S(net52261), .Z(Y[4]) );
  MUX2_X1 U48 ( .A(A[6]), .B(B[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U49 ( .A(A[9]), .B(B[9]), .S(net52635), .Z(Y[9]) );
  MUX2_X1 U50 ( .A(A[10]), .B(B[10]), .S(net52635), .Z(Y[10]) );
  MUX2_X1 U51 ( .A(A[11]), .B(B[11]), .S(net47408), .Z(Y[11]) );
  MUX2_X1 U52 ( .A(A[17]), .B(B[17]), .S(net52945), .Z(Y[17]) );
  MUX2_X1 U53 ( .A(A[20]), .B(B[20]), .S(n3), .Z(Y[20]) );
  MUX2_X1 U54 ( .A(A[22]), .B(B[22]), .S(n3), .Z(Y[22]) );
  MUX2_X1 U55 ( .A(A[23]), .B(B[23]), .S(net52463), .Z(Y[23]) );
  MUX2_X1 U56 ( .A(A[25]), .B(B[25]), .S(net52463), .Z(Y[25]) );
  MUX2_X1 U57 ( .A(A[26]), .B(B[26]), .S(net52463), .Z(Y[26]) );
  MUX2_X1 U58 ( .A(A[27]), .B(B[27]), .S(n1), .Z(Y[27]) );
  MUX2_X1 U59 ( .A(A[28]), .B(B[28]), .S(net52463), .Z(Y[28]) );
  MUX2_X1 U60 ( .A(A[31]), .B(B[31]), .S(net52261), .Z(Y[31]) );
endmodule


module MUX21_GENERIC_NBIT32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22;

  BUF_X1 U1 ( .A(n16), .Z(n9) );
  MUX2_X1 U2 ( .A(A[29]), .B(B[29]), .S(n10), .Z(Y[29]) );
  MUX2_X1 U3 ( .A(A[26]), .B(B[26]), .S(n12), .Z(Y[26]) );
  INV_X1 U4 ( .A(n14), .ZN(n1) );
  INV_X2 U5 ( .A(n19), .ZN(Y[16]) );
  INV_X1 U6 ( .A(n21), .ZN(Y[18]) );
  INV_X1 U7 ( .A(n18), .ZN(Y[9]) );
  MUX2_X2 U8 ( .A(A[10]), .B(B[10]), .S(n14), .Z(Y[10]) );
  CLKBUF_X1 U9 ( .A(n13), .Z(n12) );
  CLKBUF_X2 U10 ( .A(n13), .Z(n11) );
  MUX2_X1 U11 ( .A(A[25]), .B(B[25]), .S(n12), .Z(Y[25]) );
  NAND2_X1 U12 ( .A1(n2), .A2(n3), .ZN(Y[4]) );
  OR2_X1 U13 ( .A1(n13), .A2(n4), .ZN(n2) );
  NAND2_X1 U14 ( .A1(n13), .A2(B[4]), .ZN(n3) );
  MUX2_X1 U15 ( .A(B[8]), .B(A[8]), .S(n16), .Z(Y[8]) );
  MUX2_X2 U16 ( .A(A[23]), .B(B[23]), .S(n11), .Z(Y[23]) );
  INV_X1 U17 ( .A(A[4]), .ZN(n4) );
  INV_X1 U18 ( .A(SEL), .ZN(n16) );
  NAND2_X1 U19 ( .A1(B[19]), .A2(n15), .ZN(n6) );
  NAND2_X1 U20 ( .A1(A[19]), .A2(n9), .ZN(n7) );
  NAND2_X2 U21 ( .A1(n6), .A2(n7), .ZN(Y[19]) );
  MUX2_X2 U22 ( .A(A[24]), .B(B[24]), .S(n11), .Z(Y[24]) );
  MUX2_X2 U23 ( .A(A[20]), .B(B[20]), .S(n11), .Z(Y[20]) );
  INV_X1 U24 ( .A(n16), .ZN(n15) );
  MUX2_X2 U25 ( .A(A[22]), .B(B[22]), .S(n11), .Z(Y[22]) );
  MUX2_X1 U26 ( .A(B[15]), .B(A[15]), .S(n9), .Z(Y[15]) );
  MUX2_X2 U27 ( .A(A[27]), .B(B[27]), .S(n12), .Z(Y[27]) );
  INV_X1 U28 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U29 ( .A(n16), .ZN(n10) );
  MUX2_X2 U30 ( .A(A[21]), .B(B[21]), .S(n11), .Z(Y[21]) );
  CLKBUF_X3 U31 ( .A(SEL), .Z(n13) );
  INV_X1 U32 ( .A(n16), .ZN(n14) );
  MUX2_X1 U33 ( .A(A[0]), .B(B[0]), .S(n15), .Z(Y[0]) );
  MUX2_X1 U34 ( .A(A[1]), .B(B[1]), .S(n13), .Z(Y[1]) );
  MUX2_X1 U35 ( .A(A[2]), .B(B[2]), .S(n13), .Z(Y[2]) );
  AOI22_X1 U36 ( .A1(A[3]), .A2(n16), .B1(n13), .B2(B[3]), .ZN(n17) );
  MUX2_X1 U37 ( .A(A[5]), .B(B[5]), .S(n13), .Z(Y[5]) );
  MUX2_X1 U38 ( .A(A[6]), .B(B[6]), .S(n13), .Z(Y[6]) );
  MUX2_X1 U39 ( .A(A[7]), .B(B[7]), .S(n13), .Z(Y[7]) );
  AOI22_X1 U40 ( .A1(A[9]), .A2(n1), .B1(B[9]), .B2(n15), .ZN(n18) );
  MUX2_X1 U41 ( .A(A[11]), .B(B[11]), .S(n13), .Z(Y[11]) );
  MUX2_X1 U42 ( .A(A[12]), .B(B[12]), .S(n13), .Z(Y[12]) );
  MUX2_X1 U43 ( .A(A[13]), .B(B[13]), .S(n10), .Z(Y[13]) );
  MUX2_X1 U44 ( .A(A[14]), .B(B[14]), .S(n14), .Z(Y[14]) );
  AOI22_X1 U45 ( .A1(B[16]), .A2(n10), .B1(A[16]), .B2(n9), .ZN(n19) );
  AOI22_X1 U46 ( .A1(B[17]), .A2(n15), .B1(A[17]), .B2(n9), .ZN(n20) );
  INV_X1 U47 ( .A(n20), .ZN(Y[17]) );
  AOI22_X1 U48 ( .A1(B[18]), .A2(n15), .B1(A[18]), .B2(n9), .ZN(n21) );
  MUX2_X1 U49 ( .A(A[28]), .B(B[28]), .S(n11), .Z(Y[28]) );
  AOI22_X1 U50 ( .A1(B[30]), .A2(n10), .B1(A[30]), .B2(n9), .ZN(n22) );
  INV_X1 U51 ( .A(n22), .ZN(Y[30]) );
  MUX2_X1 U52 ( .A(A[31]), .B(B[31]), .S(n11), .Z(Y[31]) );
endmodule


module MUX21_GENERIC_NBIT32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  BUF_X2 U1 ( .A(SEL), .Z(n1) );
  BUF_X2 U2 ( .A(SEL), .Z(n2) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
  MUX2_X1 U4 ( .A(A[0]), .B(B[0]), .S(n1), .Z(Y[0]) );
  MUX2_X1 U5 ( .A(A[1]), .B(B[1]), .S(n1), .Z(Y[1]) );
  MUX2_X1 U6 ( .A(A[2]), .B(B[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U7 ( .A(A[3]), .B(B[3]), .S(n1), .Z(Y[3]) );
  MUX2_X1 U8 ( .A(A[4]), .B(B[4]), .S(n1), .Z(Y[4]) );
  MUX2_X1 U9 ( .A(A[5]), .B(B[5]), .S(n1), .Z(Y[5]) );
  MUX2_X1 U10 ( .A(A[6]), .B(B[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U11 ( .A(A[7]), .B(B[7]), .S(n1), .Z(Y[7]) );
  MUX2_X1 U12 ( .A(A[8]), .B(B[8]), .S(n1), .Z(Y[8]) );
  MUX2_X1 U13 ( .A(A[9]), .B(B[9]), .S(n1), .Z(Y[9]) );
  MUX2_X1 U14 ( .A(A[10]), .B(B[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U15 ( .A(A[11]), .B(B[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U16 ( .A(A[12]), .B(B[12]), .S(n2), .Z(Y[12]) );
  MUX2_X1 U17 ( .A(A[13]), .B(B[13]), .S(n2), .Z(Y[13]) );
  MUX2_X1 U18 ( .A(A[14]), .B(B[14]), .S(n2), .Z(Y[14]) );
  MUX2_X1 U19 ( .A(A[15]), .B(B[15]), .S(n2), .Z(Y[15]) );
  MUX2_X1 U20 ( .A(A[16]), .B(B[16]), .S(n2), .Z(Y[16]) );
  MUX2_X1 U21 ( .A(A[17]), .B(B[17]), .S(n2), .Z(Y[17]) );
  MUX2_X1 U22 ( .A(A[18]), .B(B[18]), .S(n2), .Z(Y[18]) );
  MUX2_X1 U23 ( .A(A[19]), .B(B[19]), .S(n2), .Z(Y[19]) );
  MUX2_X1 U24 ( .A(A[20]), .B(B[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U25 ( .A(A[21]), .B(B[21]), .S(n2), .Z(Y[21]) );
  MUX2_X1 U26 ( .A(A[22]), .B(B[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U27 ( .A(A[23]), .B(B[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U28 ( .A(A[24]), .B(B[24]), .S(n3), .Z(Y[24]) );
  MUX2_X1 U29 ( .A(A[25]), .B(B[25]), .S(n3), .Z(Y[25]) );
  MUX2_X1 U30 ( .A(A[26]), .B(B[26]), .S(n3), .Z(Y[26]) );
  MUX2_X1 U31 ( .A(A[27]), .B(B[27]), .S(n3), .Z(Y[27]) );
  MUX2_X1 U32 ( .A(A[28]), .B(B[28]), .S(n3), .Z(Y[28]) );
  MUX2_X1 U33 ( .A(A[29]), .B(B[29]), .S(n3), .Z(Y[29]) );
  MUX2_X1 U34 ( .A(A[30]), .B(B[30]), .S(n3), .Z(Y[30]) );
  MUX2_X1 U35 ( .A(A[31]), .B(B[31]), .S(n3), .Z(Y[31]) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  BUF_X2 U1 ( .A(SEL), .Z(n1) );
  BUF_X2 U2 ( .A(SEL), .Z(n2) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
  MUX2_X1 U4 ( .A(A[0]), .B(B[0]), .S(n1), .Z(Y[0]) );
  MUX2_X1 U5 ( .A(A[1]), .B(B[1]), .S(n1), .Z(Y[1]) );
  MUX2_X1 U6 ( .A(A[2]), .B(B[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U7 ( .A(A[3]), .B(B[3]), .S(n1), .Z(Y[3]) );
  MUX2_X1 U8 ( .A(A[4]), .B(B[4]), .S(n1), .Z(Y[4]) );
  MUX2_X1 U9 ( .A(A[5]), .B(B[5]), .S(n1), .Z(Y[5]) );
  MUX2_X1 U10 ( .A(A[6]), .B(B[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U11 ( .A(A[7]), .B(B[7]), .S(n1), .Z(Y[7]) );
  MUX2_X1 U12 ( .A(A[8]), .B(B[8]), .S(n1), .Z(Y[8]) );
  MUX2_X1 U13 ( .A(A[9]), .B(B[9]), .S(n1), .Z(Y[9]) );
  MUX2_X1 U14 ( .A(A[10]), .B(B[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U15 ( .A(A[11]), .B(B[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U16 ( .A(A[12]), .B(B[12]), .S(n2), .Z(Y[12]) );
  MUX2_X1 U17 ( .A(A[13]), .B(B[13]), .S(n2), .Z(Y[13]) );
  MUX2_X1 U18 ( .A(A[14]), .B(B[14]), .S(n2), .Z(Y[14]) );
  MUX2_X1 U19 ( .A(A[15]), .B(B[15]), .S(n2), .Z(Y[15]) );
  MUX2_X1 U20 ( .A(A[16]), .B(B[16]), .S(n2), .Z(Y[16]) );
  MUX2_X1 U21 ( .A(A[17]), .B(B[17]), .S(n2), .Z(Y[17]) );
  MUX2_X1 U22 ( .A(A[18]), .B(B[18]), .S(n2), .Z(Y[18]) );
  MUX2_X1 U23 ( .A(A[19]), .B(B[19]), .S(n2), .Z(Y[19]) );
  MUX2_X1 U24 ( .A(A[20]), .B(B[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U25 ( .A(A[21]), .B(B[21]), .S(n2), .Z(Y[21]) );
  MUX2_X1 U26 ( .A(A[22]), .B(B[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U27 ( .A(A[23]), .B(B[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U28 ( .A(A[24]), .B(B[24]), .S(n3), .Z(Y[24]) );
  MUX2_X1 U29 ( .A(A[25]), .B(B[25]), .S(n3), .Z(Y[25]) );
  MUX2_X1 U30 ( .A(A[26]), .B(B[26]), .S(n3), .Z(Y[26]) );
  MUX2_X1 U31 ( .A(A[27]), .B(B[27]), .S(n3), .Z(Y[27]) );
  MUX2_X1 U32 ( .A(A[28]), .B(B[28]), .S(n3), .Z(Y[28]) );
  MUX2_X1 U33 ( .A(A[29]), .B(B[29]), .S(n3), .Z(Y[29]) );
  MUX2_X1 U34 ( .A(A[30]), .B(B[30]), .S(n3), .Z(Y[30]) );
  MUX2_X1 U35 ( .A(A[31]), .B(B[31]), .S(n3), .Z(Y[31]) );
endmodule


module MUX21_GENERIC_NBIT5_1 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(A[0]), .B(B[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(A[1]), .B(B[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(A[2]), .B(B[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(A[3]), .B(B[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U5 ( .A(A[4]), .B(B[4]), .S(SEL), .Z(Y[4]) );
endmodule


module ADDER_N32_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2_X2 U2 ( .A1(A[2]), .A2(A[3]), .ZN(n1) );
  AND4_X1 U3 ( .A1(A[11]), .A2(n13), .A3(n14), .A4(A[8]), .ZN(n2) );
  NAND4_X1 U4 ( .A1(A[11]), .A2(n13), .A3(n14), .A4(A[8]), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n23), .A2(n2), .ZN(n4) );
  BUF_X2 U6 ( .A(A[9]), .Z(n14) );
  BUF_X2 U7 ( .A(A[10]), .Z(n13) );
  AND2_X1 U8 ( .A1(n19), .A2(n5), .ZN(n35) );
  AND2_X1 U9 ( .A1(n37), .A2(n7), .ZN(n5) );
  INV_X1 U10 ( .A(n54), .ZN(n64) );
  AND4_X1 U11 ( .A1(n43), .A2(n44), .A3(n45), .A4(A[27]), .ZN(n6) );
  AND2_X1 U12 ( .A1(n6), .A2(n40), .ZN(n7) );
  XNOR2_X1 U13 ( .A(n63), .B(n61), .ZN(SUM[22]) );
  XNOR2_X1 U14 ( .A(n48), .B(n22), .ZN(SUM[26]) );
  NOR2_X1 U15 ( .A1(n87), .A2(n27), .ZN(n8) );
  AND2_X1 U16 ( .A1(n19), .A2(n7), .ZN(n39) );
  AND2_X1 U17 ( .A1(n19), .A2(n43), .ZN(n49) );
  INV_X1 U18 ( .A(n17), .ZN(n9) );
  AND2_X1 U19 ( .A1(n19), .A2(n6), .ZN(n42) );
  XNOR2_X1 U20 ( .A(n25), .B(n70), .ZN(SUM[19]) );
  AND2_X1 U21 ( .A1(n24), .A2(n10), .ZN(n60) );
  AND2_X1 U22 ( .A1(n56), .A2(n58), .ZN(n10) );
  XNOR2_X1 U23 ( .A(n62), .B(n60), .ZN(SUM[23]) );
  XNOR2_X1 U24 ( .A(n11), .B(n47), .ZN(SUM[27]) );
  AND2_X1 U25 ( .A1(n45), .A2(n22), .ZN(n11) );
  CLKBUF_X1 U26 ( .A(n14), .Z(n12) );
  AND4_X2 U27 ( .A1(A[4]), .A2(A[5]), .A3(A[6]), .A4(A[7]), .ZN(n23) );
  NOR2_X1 U28 ( .A1(n67), .A2(n15), .ZN(n71) );
  OR2_X1 U29 ( .A1(n73), .A2(n74), .ZN(n15) );
  XNOR2_X1 U30 ( .A(n16), .B(n34), .ZN(SUM[31]) );
  AND2_X1 U31 ( .A1(n35), .A2(n36), .ZN(n16) );
  NOR2_X1 U32 ( .A1(n75), .A2(n76), .ZN(n17) );
  NOR2_X1 U33 ( .A1(n4), .A2(n76), .ZN(n18) );
  NOR2_X1 U34 ( .A1(n75), .A2(n76), .ZN(n51) );
  AND2_X2 U35 ( .A1(n51), .A2(n52), .ZN(n19) );
  NOR2_X1 U36 ( .A1(n67), .A2(n54), .ZN(n66) );
  NOR2_X1 U37 ( .A1(n83), .A2(n86), .ZN(n82) );
  AND2_X1 U38 ( .A1(n23), .A2(n1), .ZN(n20) );
  NAND2_X1 U39 ( .A1(n23), .A2(n1), .ZN(n87) );
  OR2_X1 U40 ( .A1(n87), .A2(n3), .ZN(n21) );
  NAND2_X1 U41 ( .A1(n23), .A2(n2), .ZN(n75) );
  NOR2_X1 U42 ( .A1(n9), .A2(n73), .ZN(n72) );
  AND3_X1 U43 ( .A1(n19), .A2(n43), .A3(n44), .ZN(n22) );
  NOR2_X1 U44 ( .A1(n53), .A2(n54), .ZN(n52) );
  NAND4_X1 U45 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(n53) );
  AND2_X1 U46 ( .A1(n24), .A2(n56), .ZN(n61) );
  AND3_X1 U47 ( .A1(n55), .A2(n64), .A3(n18), .ZN(n24) );
  AND2_X1 U48 ( .A1(n71), .A2(A[18]), .ZN(n25) );
  NAND4_X1 U49 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n68), .ZN(n54) );
  NOR2_X1 U50 ( .A1(n87), .A2(n27), .ZN(n26) );
  OR2_X1 U51 ( .A1(n77), .A2(n3), .ZN(n27) );
  AND2_X1 U52 ( .A1(n1), .A2(A[4]), .ZN(n28) );
  AND2_X1 U53 ( .A1(n80), .A2(n26), .ZN(n29) );
  AND2_X1 U54 ( .A1(n30), .A2(n14), .ZN(n89) );
  AND2_X1 U55 ( .A1(n28), .A2(A[5]), .ZN(n33) );
  AND2_X1 U56 ( .A1(n20), .A2(A[8]), .ZN(n30) );
  AND2_X1 U57 ( .A1(A[6]), .A2(n33), .ZN(n31) );
  AND2_X1 U58 ( .A1(n13), .A2(n89), .ZN(n32) );
  INV_X1 U59 ( .A(A[12]), .ZN(n77) );
  INV_X1 U60 ( .A(n59), .ZN(n43) );
  INV_X1 U61 ( .A(A[24]), .ZN(n59) );
  INV_X1 U62 ( .A(n48), .ZN(n45) );
  INV_X1 U63 ( .A(A[26]), .ZN(n48) );
  INV_X1 U64 ( .A(n63), .ZN(n58) );
  INV_X1 U65 ( .A(A[22]), .ZN(n63) );
  INV_X1 U66 ( .A(n65), .ZN(n56) );
  INV_X1 U67 ( .A(A[21]), .ZN(n65) );
  INV_X1 U68 ( .A(A[17]), .ZN(n74) );
  INV_X1 U69 ( .A(n50), .ZN(n44) );
  INV_X1 U70 ( .A(A[25]), .ZN(n50) );
  INV_X1 U71 ( .A(n88), .ZN(n80) );
  INV_X1 U72 ( .A(A[13]), .ZN(n88) );
  INV_X1 U73 ( .A(n69), .ZN(n55) );
  INV_X1 U74 ( .A(A[20]), .ZN(n69) );
  INV_X1 U75 ( .A(n70), .ZN(n68) );
  INV_X1 U76 ( .A(A[19]), .ZN(n70) );
  INV_X1 U77 ( .A(n46), .ZN(n40) );
  INV_X1 U78 ( .A(A[28]), .ZN(n46) );
  INV_X1 U79 ( .A(n38), .ZN(n36) );
  INV_X1 U80 ( .A(A[30]), .ZN(n38) );
  INV_X1 U81 ( .A(n86), .ZN(n84) );
  INV_X1 U82 ( .A(A[14]), .ZN(n86) );
  INV_X1 U83 ( .A(n85), .ZN(n81) );
  INV_X1 U84 ( .A(A[15]), .ZN(n85) );
  INV_X1 U85 ( .A(n41), .ZN(n37) );
  INV_X1 U86 ( .A(A[29]), .ZN(n41) );
  INV_X1 U87 ( .A(n62), .ZN(n57) );
  INV_X1 U88 ( .A(A[23]), .ZN(n62) );
  INV_X1 U89 ( .A(A[31]), .ZN(n34) );
  XOR2_X1 U90 ( .A(n36), .B(n35), .Z(SUM[30]) );
  XOR2_X1 U91 ( .A(n40), .B(n42), .Z(SUM[28]) );
  XOR2_X1 U92 ( .A(n44), .B(n49), .Z(SUM[25]) );
  XOR2_X1 U93 ( .A(n37), .B(n39), .Z(SUM[29]) );
  XOR2_X1 U94 ( .A(A[16]), .B(n17), .Z(SUM[16]) );
  XOR2_X1 U95 ( .A(n13), .B(n89), .Z(SUM[10]) );
  XOR2_X1 U96 ( .A(n24), .B(n56), .Z(SUM[21]) );
  XOR2_X1 U97 ( .A(A[2]), .B(A[3]), .Z(SUM[3]) );
  XOR2_X1 U98 ( .A(A[8]), .B(n20), .Z(SUM[8]) );
  XOR2_X1 U99 ( .A(A[4]), .B(n1), .Z(SUM[4]) );
  XOR2_X1 U100 ( .A(n43), .B(n19), .Z(SUM[24]) );
  XOR2_X1 U101 ( .A(A[6]), .B(n33), .Z(SUM[6]) );
  XOR2_X1 U102 ( .A(n84), .B(n29), .Z(SUM[14]) );
  INV_X1 U103 ( .A(A[2]), .ZN(SUM[2]) );
  XOR2_X1 U104 ( .A(n81), .B(n82), .Z(SUM[15]) );
  XOR2_X1 U105 ( .A(A[17]), .B(n72), .Z(SUM[17]) );
  XOR2_X1 U106 ( .A(n55), .B(n66), .Z(SUM[20]) );
  XOR2_X1 U107 ( .A(A[11]), .B(n32), .Z(SUM[11]) );
  XOR2_X1 U108 ( .A(A[18]), .B(n71), .Z(SUM[18]) );
  XOR2_X1 U109 ( .A(A[7]), .B(n31), .Z(SUM[7]) );
  XOR2_X1 U110 ( .A(n30), .B(n12), .Z(SUM[9]) );
  XOR2_X1 U111 ( .A(n80), .B(n8), .Z(SUM[13]) );
  XOR2_X1 U112 ( .A(n21), .B(n77), .Z(SUM[12]) );
  XOR2_X1 U113 ( .A(A[5]), .B(n28), .Z(SUM[5]) );
  INV_X1 U114 ( .A(A[27]), .ZN(n47) );
  INV_X1 U115 ( .A(A[16]), .ZN(n73) );
  INV_X1 U116 ( .A(n18), .ZN(n67) );
  NAND3_X1 U117 ( .A1(n1), .A2(n78), .A3(n79), .ZN(n76) );
  NOR2_X1 U118 ( .A1(n88), .A2(n77), .ZN(n79) );
  NOR2_X1 U119 ( .A1(n85), .A2(n86), .ZN(n78) );
  INV_X1 U120 ( .A(n29), .ZN(n83) );
endmodule


module ADDER_N32 ( CURR_ADDR, NEXT_ADDR );
  input [31:0] CURR_ADDR;
  output [31:0] NEXT_ADDR;


  ADDER_N32_DW01_add_2 add_26 ( .A(CURR_ADDR), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(NEXT_ADDR) );
endmodule


module REGISTER_FILE_NBIT32_NREG32 ( CLK, RST, EN, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST, EN, RD1, RD2, WR;
  wire   n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462;

  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n3614), .CK(CLK), .QN(n2168) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n3613), .CK(CLK), .QN(n2126) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n3612), .CK(CLK), .QN(n2090) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n3611), .CK(CLK), .QN(n2054) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n3610), .CK(CLK), .QN(n2018) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n3609), .CK(CLK), .QN(n1982) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n3608), .CK(CLK), .QN(n1946) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n3607), .CK(CLK), .QN(n1910) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n3606), .CK(CLK), .QN(n1874) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n3605), .CK(CLK), .QN(n1838) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n3604), .CK(CLK), .QN(n1802) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n3603), .CK(CLK), .QN(n1766) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n3602), .CK(CLK), .QN(n1730) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n3601), .CK(CLK), .QN(n1694) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n3600), .CK(CLK), .QN(n1658) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n3599), .CK(CLK), .QN(n1622) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n3598), .CK(CLK), .QN(n1586) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n3597), .CK(CLK), .QN(n1550) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n3596), .CK(CLK), .QN(n1514) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n3595), .CK(CLK), .QN(n1478) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n3594), .CK(CLK), .QN(n1442) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n3593), .CK(CLK), .QN(n1406) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n3592), .CK(CLK), .QN(n1370) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n3591), .CK(CLK), .QN(n1334) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n3590), .CK(CLK), .QN(n1298) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n3589), .CK(CLK), .QN(n1262) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n3588), .CK(CLK), .QN(n1226) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n3587), .CK(CLK), .QN(n1190) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n3586), .CK(CLK), .QN(n1154) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n3585), .CK(CLK), .QN(n1118) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n3584), .CK(CLK), .QN(n1082) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n3583), .CK(CLK), .QN(n1044) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n3582), .CK(CLK), .QN(n2170) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n3581), .CK(CLK), .QN(n2127) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n3580), .CK(CLK), .QN(n2091) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n3579), .CK(CLK), .QN(n2055) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n3578), .CK(CLK), .QN(n2019) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n3577), .CK(CLK), .QN(n1983) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n3576), .CK(CLK), .QN(n1947) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n3575), .CK(CLK), .QN(n1911) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n3574), .CK(CLK), .QN(n1875) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n3573), .CK(CLK), .QN(n1839) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n3572), .CK(CLK), .QN(n1803) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n3571), .CK(CLK), .QN(n1767) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n3570), .CK(CLK), .QN(n1731) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n3569), .CK(CLK), .QN(n1695) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n3568), .CK(CLK), .QN(n1659) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n3567), .CK(CLK), .QN(n1623) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n3566), .CK(CLK), .QN(n1587) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n3565), .CK(CLK), .QN(n1551) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n3564), .CK(CLK), .QN(n1515) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n3563), .CK(CLK), .QN(n1479) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n3562), .CK(CLK), .QN(n1443) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n3561), .CK(CLK), .QN(n1407) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n3560), .CK(CLK), .QN(n1371) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n3559), .CK(CLK), .QN(n1335) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n3558), .CK(CLK), .QN(n1299) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n3557), .CK(CLK), .QN(n1263) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n3556), .CK(CLK), .QN(n1227) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n3555), .CK(CLK), .QN(n1191) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n3554), .CK(CLK), .QN(n1155) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n3553), .CK(CLK), .QN(n1119) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n3552), .CK(CLK), .QN(n1083) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n3551), .CK(CLK), .QN(n1045) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n3550), .CK(CLK), .Q(n4358) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n3549), .CK(CLK), .Q(n4355) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n3548), .CK(CLK), .Q(n4353) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n3547), .CK(CLK), .Q(n4351) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n3546), .CK(CLK), .Q(n4349) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n3545), .CK(CLK), .Q(n4347) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n3544), .CK(CLK), .Q(n4345) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n3543), .CK(CLK), .Q(n4343) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n3542), .CK(CLK), .Q(n4341) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n3541), .CK(CLK), .Q(n4339) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n3540), .CK(CLK), .Q(n4337) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n3539), .CK(CLK), .Q(n4335) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n3538), .CK(CLK), .Q(n4333) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n3537), .CK(CLK), .Q(n4331) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n3536), .CK(CLK), .Q(n4329) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n3535), .CK(CLK), .Q(n4327) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n3534), .CK(CLK), .Q(n4325) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n3533), .CK(CLK), .Q(n4323) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n3532), .CK(CLK), .Q(n4321) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n3531), .CK(CLK), .Q(n4319) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n3530), .CK(CLK), .Q(n4317) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n3529), .CK(CLK), .Q(n4315) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n3528), .CK(CLK), .Q(n4313) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n3527), .CK(CLK), .Q(n4311) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n3526), .CK(CLK), .Q(n4309) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n3525), .CK(CLK), .Q(n4307) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n3524), .CK(CLK), .Q(n4305) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n3523), .CK(CLK), .Q(n4303) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n3522), .CK(CLK), .Q(n4301) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n3521), .CK(CLK), .Q(n4299) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n3520), .CK(CLK), .Q(n4297) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n3519), .CK(CLK), .Q(n4295) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n3518), .CK(CLK), .Q(n4292) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n3517), .CK(CLK), .Q(n4290) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n3516), .CK(CLK), .Q(n4289) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n3515), .CK(CLK), .Q(n4288) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n3514), .CK(CLK), .Q(n4287) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n3513), .CK(CLK), .Q(n4286) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n3512), .CK(CLK), .Q(n4285) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n3511), .CK(CLK), .Q(n4284) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n3510), .CK(CLK), .Q(n4283) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n3509), .CK(CLK), .Q(n4282) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n3508), .CK(CLK), .Q(n4281) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n3507), .CK(CLK), .Q(n4280) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n3506), .CK(CLK), .Q(n4279) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n3505), .CK(CLK), .Q(n4278) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n3504), .CK(CLK), .Q(n4277) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n3503), .CK(CLK), .Q(n4276) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n3502), .CK(CLK), .Q(n4275) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n3501), .CK(CLK), .Q(n4274) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n3500), .CK(CLK), .Q(n4273) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n3499), .CK(CLK), .Q(n4272) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n3498), .CK(CLK), .Q(n4271) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n3497), .CK(CLK), .Q(n4270) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n3496), .CK(CLK), .Q(n4269) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n3495), .CK(CLK), .Q(n4268) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n3494), .CK(CLK), .Q(n4267) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n3493), .CK(CLK), .Q(n4266) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n3492), .CK(CLK), .Q(n4265) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n3491), .CK(CLK), .Q(n4264) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n3490), .CK(CLK), .Q(n4263) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n3489), .CK(CLK), .Q(n4262) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n3488), .CK(CLK), .Q(n4261) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n3487), .CK(CLK), .Q(n4260) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n3486), .CK(CLK), .QN(n2163) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n3485), .CK(CLK), .QN(n2123) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n3484), .CK(CLK), .QN(n2087) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n3483), .CK(CLK), .QN(n2051) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n3482), .CK(CLK), .QN(n2015) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n3481), .CK(CLK), .QN(n1979) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n3480), .CK(CLK), .QN(n1943) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n3479), .CK(CLK), .QN(n1907) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n3478), .CK(CLK), .QN(n1871) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n3477), .CK(CLK), .QN(n1835) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n3476), .CK(CLK), .QN(n1799) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n3475), .CK(CLK), .QN(n1763) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n3474), .CK(CLK), .QN(n1727) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n3473), .CK(CLK), .QN(n1691) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n3472), .CK(CLK), .QN(n1655) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n3471), .CK(CLK), .QN(n1619) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n3470), .CK(CLK), .QN(n1583) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n3469), .CK(CLK), .QN(n1547) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n3468), .CK(CLK), .QN(n1511) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n3467), .CK(CLK), .QN(n1475) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n3466), .CK(CLK), .QN(n1439) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n3465), .CK(CLK), .QN(n1403) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n3464), .CK(CLK), .QN(n1367) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n3463), .CK(CLK), .QN(n1331) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n3462), .CK(CLK), .QN(n1295) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n3461), .CK(CLK), .QN(n1259) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n3460), .CK(CLK), .QN(n1223) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n3459), .CK(CLK), .QN(n1187) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n3458), .CK(CLK), .QN(n1151) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n3457), .CK(CLK), .QN(n1115) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n3456), .CK(CLK), .QN(n1079) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n3455), .CK(CLK), .QN(n1041) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n3454), .CK(CLK), .QN(n2165) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n3453), .CK(CLK), .QN(n2124) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n3452), .CK(CLK), .QN(n2088) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n3451), .CK(CLK), .QN(n2052) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n3450), .CK(CLK), .QN(n2016) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n3449), .CK(CLK), .QN(n1980) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n3448), .CK(CLK), .QN(n1944) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n3447), .CK(CLK), .QN(n1908) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n3446), .CK(CLK), .QN(n1872) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n3445), .CK(CLK), .QN(n1836) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n3444), .CK(CLK), .QN(n1800) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n3443), .CK(CLK), .QN(n1764) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n3442), .CK(CLK), .QN(n1728) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n3441), .CK(CLK), .QN(n1692) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n3440), .CK(CLK), .QN(n1656) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n3439), .CK(CLK), .QN(n1620) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n3438), .CK(CLK), .QN(n1584) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n3437), .CK(CLK), .QN(n1548) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n3436), .CK(CLK), .QN(n1512) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n3435), .CK(CLK), .QN(n1476) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n3434), .CK(CLK), .QN(n1440) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n3433), .CK(CLK), .QN(n1404) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n3432), .CK(CLK), .QN(n1368) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n3431), .CK(CLK), .QN(n1332) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n3430), .CK(CLK), .QN(n1296) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n3429), .CK(CLK), .QN(n1260) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n3428), .CK(CLK), .QN(n1224) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n3427), .CK(CLK), .QN(n1188) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n3426), .CK(CLK), .QN(n1152) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n3425), .CK(CLK), .QN(n1116) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n3424), .CK(CLK), .QN(n1080) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n3423), .CK(CLK), .QN(n1042) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n3422), .CK(CLK), .Q(n4187) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n3421), .CK(CLK), .Q(n4185) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n3420), .CK(CLK), .Q(n4184) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n3419), .CK(CLK), .Q(n4183) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n3418), .CK(CLK), .Q(n4182) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n3417), .CK(CLK), .Q(n4181) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n3416), .CK(CLK), .Q(n4180) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n3415), .CK(CLK), .Q(n4179) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n3414), .CK(CLK), .Q(n4178) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n3413), .CK(CLK), .Q(n4177) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n3412), .CK(CLK), .Q(n4176) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n3411), .CK(CLK), .Q(n4175) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n3410), .CK(CLK), .Q(n4174) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n3409), .CK(CLK), .Q(n4173) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n3408), .CK(CLK), .Q(n4172) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n3407), .CK(CLK), .Q(n4171) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n3406), .CK(CLK), .Q(n4170) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n3405), .CK(CLK), .Q(n4169) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n3404), .CK(CLK), .Q(n4168) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n3403), .CK(CLK), .Q(n4167) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n3402), .CK(CLK), .Q(n4166) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n3401), .CK(CLK), .Q(n4165) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n3400), .CK(CLK), .Q(n4164) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n3399), .CK(CLK), .Q(n4163) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n3398), .CK(CLK), .Q(n4162) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n3397), .CK(CLK), .Q(n4161) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n3396), .CK(CLK), .Q(n4160) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n3395), .CK(CLK), .Q(n4159) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n3394), .CK(CLK), .Q(n4158) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n3393), .CK(CLK), .Q(n4157) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n3392), .CK(CLK), .Q(n4156) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n3391), .CK(CLK), .Q(n4155) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n3390), .CK(CLK), .Q(n4152) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n3389), .CK(CLK), .Q(n4150) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n3388), .CK(CLK), .Q(n4149) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n3387), .CK(CLK), .Q(n4148) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n3386), .CK(CLK), .Q(n4147) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n3385), .CK(CLK), .Q(n4146) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n3384), .CK(CLK), .Q(n4145) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n3383), .CK(CLK), .Q(n4144) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n3382), .CK(CLK), .Q(n4143) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n3381), .CK(CLK), .Q(n4142) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n3380), .CK(CLK), .Q(n4141) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n3379), .CK(CLK), .Q(n4140) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n3378), .CK(CLK), .Q(n4139) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n3377), .CK(CLK), .Q(n4138) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n3376), .CK(CLK), .Q(n4137) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n3375), .CK(CLK), .Q(n4136) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n3374), .CK(CLK), .Q(n4135) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n3373), .CK(CLK), .Q(n4134) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n3372), .CK(CLK), .Q(n4133) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n3371), .CK(CLK), .Q(n4132) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n3370), .CK(CLK), .Q(n4131) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n3369), .CK(CLK), .Q(n4130) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n3368), .CK(CLK), .Q(n4129) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n3367), .CK(CLK), .Q(n4128) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n3366), .CK(CLK), .Q(n4127) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n3365), .CK(CLK), .Q(n4126) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n3364), .CK(CLK), .Q(n4125) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n3363), .CK(CLK), .Q(n4124) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n3362), .CK(CLK), .Q(n4123) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n3361), .CK(CLK), .Q(n4122) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n3360), .CK(CLK), .Q(n4121) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n3359), .CK(CLK), .Q(n4120) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n3358), .CK(CLK), .QN(n2158) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n3357), .CK(CLK), .QN(n2120) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n3356), .CK(CLK), .QN(n2084) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n3355), .CK(CLK), .QN(n2048) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n3354), .CK(CLK), .QN(n2012) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n3353), .CK(CLK), .QN(n1976) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n3352), .CK(CLK), .QN(n1940) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n3351), .CK(CLK), .QN(n1904) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n3350), .CK(CLK), .QN(n1868) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n3349), .CK(CLK), .QN(n1832) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n3348), .CK(CLK), .QN(n1796) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n3347), .CK(CLK), .QN(n1760) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n3346), .CK(CLK), .QN(n1724) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n3345), .CK(CLK), .QN(n1688) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n3344), .CK(CLK), .QN(n1652) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n3343), .CK(CLK), .QN(n1616) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n3342), .CK(CLK), .QN(n1580) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n3341), .CK(CLK), .QN(n1544) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n3340), .CK(CLK), .QN(n1508) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n3339), .CK(CLK), .QN(n1472) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n3338), .CK(CLK), .QN(n1436) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n3337), .CK(CLK), .QN(n1400) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n3336), .CK(CLK), .QN(n1364) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n3335), .CK(CLK), .QN(n1328) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n3334), .CK(CLK), .QN(n1292) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n3333), .CK(CLK), .QN(n1256) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n3332), .CK(CLK), .QN(n1220) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n3331), .CK(CLK), .QN(n1184) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n3330), .CK(CLK), .QN(n1148) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n3329), .CK(CLK), .QN(n1112) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n3328), .CK(CLK), .QN(n1076) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n3327), .CK(CLK), .QN(n1037) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n3326), .CK(CLK), .QN(n2160) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n3325), .CK(CLK), .QN(n2121) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n3324), .CK(CLK), .QN(n2085) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n3323), .CK(CLK), .QN(n2049) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n3322), .CK(CLK), .QN(n2013) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n3321), .CK(CLK), .QN(n1977) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n3320), .CK(CLK), .QN(n1941) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n3319), .CK(CLK), .QN(n1905) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n3318), .CK(CLK), .QN(n1869) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n3317), .CK(CLK), .QN(n1833) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n3316), .CK(CLK), .QN(n1797) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n3315), .CK(CLK), .QN(n1761) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n3314), .CK(CLK), .QN(n1725) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n3313), .CK(CLK), .QN(n1689) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n3312), .CK(CLK), .QN(n1653) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n3311), .CK(CLK), .QN(n1617) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n3310), .CK(CLK), .QN(n1581) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n3309), .CK(CLK), .QN(n1545) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n3308), .CK(CLK), .QN(n1509) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n3307), .CK(CLK), .QN(n1473) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n3306), .CK(CLK), .QN(n1437) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n3305), .CK(CLK), .QN(n1401) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n3304), .CK(CLK), .QN(n1365) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n3303), .CK(CLK), .QN(n1329) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n3302), .CK(CLK), .QN(n1293) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n3301), .CK(CLK), .QN(n1257) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n3300), .CK(CLK), .QN(n1221) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n3299), .CK(CLK), .QN(n1185) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n3298), .CK(CLK), .QN(n1149) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n3297), .CK(CLK), .QN(n1113) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n3296), .CK(CLK), .QN(n1077) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n3295), .CK(CLK), .QN(n1038) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n3294), .CK(CLK), .Q(n4046) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n3293), .CK(CLK), .Q(n4044) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n3292), .CK(CLK), .Q(n4043) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n3291), .CK(CLK), .Q(n4042) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n3290), .CK(CLK), .Q(n4041) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n3289), .CK(CLK), .Q(n4040) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n3288), .CK(CLK), .Q(n4039) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n3287), .CK(CLK), .Q(n4038) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n3286), .CK(CLK), .Q(n4037) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n3285), .CK(CLK), .Q(n4036) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n3284), .CK(CLK), .Q(n4035) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n3283), .CK(CLK), .Q(n4034) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n3282), .CK(CLK), .Q(n4033) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n3281), .CK(CLK), .Q(n4032) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n3280), .CK(CLK), .Q(n4031) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n3279), .CK(CLK), .Q(n4030) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n3278), .CK(CLK), .Q(n4029) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n3277), .CK(CLK), .Q(n4028) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n3276), .CK(CLK), .Q(n4027) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n3275), .CK(CLK), .Q(n4026) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n3274), .CK(CLK), .Q(n4025) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n3273), .CK(CLK), .Q(n4024) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n3272), .CK(CLK), .Q(n4023) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n3271), .CK(CLK), .Q(n4022) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n3270), .CK(CLK), .Q(n4021) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n3269), .CK(CLK), .Q(n4020) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n3268), .CK(CLK), .Q(n4019) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n3267), .CK(CLK), .Q(n4018) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n3266), .CK(CLK), .Q(n4017) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n3265), .CK(CLK), .Q(n4016) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n3264), .CK(CLK), .Q(n4015) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n3263), .CK(CLK), .Q(n4014) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n3262), .CK(CLK), .Q(n4012) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n3261), .CK(CLK), .Q(n4010) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n3260), .CK(CLK), .Q(n4009) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n3259), .CK(CLK), .Q(n4008) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n3258), .CK(CLK), .Q(n4007) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n3257), .CK(CLK), .Q(n4006) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n3256), .CK(CLK), .Q(n4005) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n3255), .CK(CLK), .Q(n4004) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n3254), .CK(CLK), .Q(n4003) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n3253), .CK(CLK), .Q(n4002) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n3252), .CK(CLK), .Q(n4001) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n3251), .CK(CLK), .Q(n4000) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n3250), .CK(CLK), .Q(n3999) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n3249), .CK(CLK), .Q(n3998) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n3248), .CK(CLK), .Q(n3997) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n3247), .CK(CLK), .Q(n3996) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n3246), .CK(CLK), .Q(n3995) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n3245), .CK(CLK), .Q(n3994) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n3244), .CK(CLK), .Q(n3993) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n3243), .CK(CLK), .Q(n3992) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n3242), .CK(CLK), .Q(n3991) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n3241), .CK(CLK), .Q(n3990) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n3240), .CK(CLK), .Q(n3989) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n3239), .CK(CLK), .Q(n3988) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n3238), .CK(CLK), .Q(n3987) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n3237), .CK(CLK), .Q(n3986) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n3236), .CK(CLK), .Q(n3985) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n3235), .CK(CLK), .Q(n3984) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n3234), .CK(CLK), .Q(n3983) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n3233), .CK(CLK), .Q(n3982) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n3232), .CK(CLK), .Q(n3981) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n3231), .CK(CLK), .Q(n3980) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n3230), .CK(CLK), .QN(n2153) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n3229), .CK(CLK), .QN(n2117) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n3228), .CK(CLK), .QN(n2081) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n3227), .CK(CLK), .QN(n2045) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n3226), .CK(CLK), .QN(n2009) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n3225), .CK(CLK), .QN(n1973) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n3224), .CK(CLK), .QN(n1937) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n3223), .CK(CLK), .QN(n1901) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n3222), .CK(CLK), .QN(n1865) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n3221), .CK(CLK), .QN(n1829) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n3220), .CK(CLK), .QN(n1793) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n3219), .CK(CLK), .QN(n1757) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n3218), .CK(CLK), .QN(n1721) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n3217), .CK(CLK), .QN(n1685) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n3216), .CK(CLK), .QN(n1649) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n3215), .CK(CLK), .QN(n1613) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n3214), .CK(CLK), .QN(n1577) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n3213), .CK(CLK), .QN(n1541) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n3212), .CK(CLK), .QN(n1505) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n3211), .CK(CLK), .QN(n1469) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n3210), .CK(CLK), .QN(n1433) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n3209), .CK(CLK), .QN(n1397) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n3208), .CK(CLK), .QN(n1361) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n3207), .CK(CLK), .QN(n1325) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n3206), .CK(CLK), .QN(n1289) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n3205), .CK(CLK), .QN(n1253) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n3204), .CK(CLK), .QN(n1217) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n3203), .CK(CLK), .QN(n1181) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n3202), .CK(CLK), .QN(n1145) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n3201), .CK(CLK), .QN(n1109) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n3200), .CK(CLK), .QN(n1073) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n3199), .CK(CLK), .QN(n1032) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n3198), .CK(CLK), .QN(n2155) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n3197), .CK(CLK), .QN(n2118) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n3196), .CK(CLK), .QN(n2082) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n3195), .CK(CLK), .QN(n2046) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n3194), .CK(CLK), .QN(n2010) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n3193), .CK(CLK), .QN(n1974) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n3192), .CK(CLK), .QN(n1938) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n3191), .CK(CLK), .QN(n1902) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n3190), .CK(CLK), .QN(n1866) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n3189), .CK(CLK), .QN(n1830) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n3188), .CK(CLK), .QN(n1794) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n3187), .CK(CLK), .QN(n1758) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n3186), .CK(CLK), .QN(n1722) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n3185), .CK(CLK), .QN(n1686) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n3184), .CK(CLK), .QN(n1650) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n3183), .CK(CLK), .QN(n1614) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n3182), .CK(CLK), .QN(n1578) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n3181), .CK(CLK), .QN(n1542) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n3180), .CK(CLK), .QN(n1506) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n3179), .CK(CLK), .QN(n1470) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n3178), .CK(CLK), .QN(n1434) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n3177), .CK(CLK), .QN(n1398) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n3176), .CK(CLK), .QN(n1362) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n3175), .CK(CLK), .QN(n1326) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n3174), .CK(CLK), .QN(n1290) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n3173), .CK(CLK), .QN(n1254) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n3172), .CK(CLK), .QN(n1218) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n3171), .CK(CLK), .QN(n1182) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n3170), .CK(CLK), .QN(n1146) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n3169), .CK(CLK), .QN(n1110) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n3168), .CK(CLK), .QN(n1074) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n3167), .CK(CLK), .QN(n1033) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n3166), .CK(CLK), .Q(n3910) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n3165), .CK(CLK), .Q(n3908) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n3164), .CK(CLK), .Q(n3907) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n3163), .CK(CLK), .Q(n3906) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n3162), .CK(CLK), .Q(n3905) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n3161), .CK(CLK), .Q(n3904) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n3160), .CK(CLK), .Q(n3903) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n3159), .CK(CLK), .Q(n3902) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n3158), .CK(CLK), .Q(n3901) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n3157), .CK(CLK), .Q(n3900) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n3156), .CK(CLK), .Q(n3899) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n3155), .CK(CLK), .Q(n3898) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n3154), .CK(CLK), .Q(n3897) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n3153), .CK(CLK), .Q(n3896) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n3152), .CK(CLK), .Q(n3895) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n3151), .CK(CLK), .Q(n3894) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n3150), .CK(CLK), .Q(n3893) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n3149), .CK(CLK), .Q(n3892) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n3148), .CK(CLK), .Q(n3891) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n3147), .CK(CLK), .Q(n3890) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n3146), .CK(CLK), .Q(n3889) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n3145), .CK(CLK), .Q(n3888) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n3144), .CK(CLK), .Q(n3887) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n3143), .CK(CLK), .Q(n3886) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n3142), .CK(CLK), .Q(n3885) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n3141), .CK(CLK), .Q(n3884) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n3140), .CK(CLK), .Q(n3883) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n3139), .CK(CLK), .Q(n3882) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n3138), .CK(CLK), .Q(n3881) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n3137), .CK(CLK), .Q(n3880) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n3136), .CK(CLK), .Q(n3879) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n3135), .CK(CLK), .Q(n3878) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n3134), .CK(CLK), .Q(n3876) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n3133), .CK(CLK), .Q(n3874) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n3132), .CK(CLK), .Q(n3873) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n3131), .CK(CLK), .Q(n3872) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n3130), .CK(CLK), .Q(n3871) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n3129), .CK(CLK), .Q(n3870) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n3128), .CK(CLK), .Q(n3869) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n3127), .CK(CLK), .Q(n3868) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n3126), .CK(CLK), .Q(n3867) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n3125), .CK(CLK), .Q(n3866) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n3124), .CK(CLK), .Q(n3865) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n3123), .CK(CLK), .Q(n3864) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n3122), .CK(CLK), .Q(n3863) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n3121), .CK(CLK), .Q(n3862) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n3120), .CK(CLK), .Q(n3861) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n3119), .CK(CLK), .Q(n3860) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n3118), .CK(CLK), .Q(n3859) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n3117), .CK(CLK), .Q(n3858) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n3116), .CK(CLK), .Q(n3857) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n3115), .CK(CLK), .Q(n3856) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n3114), .CK(CLK), .Q(n3855) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n3113), .CK(CLK), .Q(n3854) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n3112), .CK(CLK), .Q(n3853) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n3111), .CK(CLK), .Q(n3852) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n3110), .CK(CLK), .Q(n3851) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n3109), .CK(CLK), .Q(n3850) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n3108), .CK(CLK), .Q(n3849) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n3107), .CK(CLK), .Q(n3848) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n3106), .CK(CLK), .Q(n3847) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n3105), .CK(CLK), .Q(n3846) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n3104), .CK(CLK), .Q(n3845) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n3103), .CK(CLK), .Q(n3844) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n3102), .CK(CLK), .QN(n2192) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n3101), .CK(CLK), .QN(n2142) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n3100), .CK(CLK), .QN(n2106) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n3099), .CK(CLK), .QN(n2070) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n3098), .CK(CLK), .QN(n2034) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n3097), .CK(CLK), .QN(n1998) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n3096), .CK(CLK), .QN(n1962) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n3095), .CK(CLK), .QN(n1926) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n3094), .CK(CLK), .QN(n1890) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n3093), .CK(CLK), .QN(n1854) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n3092), .CK(CLK), .QN(n1818) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n3091), .CK(CLK), .QN(n1782) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n3090), .CK(CLK), .QN(n1746) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n3089), .CK(CLK), .QN(n1710) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n3088), .CK(CLK), .QN(n1674) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n3087), .CK(CLK), .QN(n1638) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n3086), .CK(CLK), .QN(n1602) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n3085), .CK(CLK), .QN(n1566) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n3084), .CK(CLK), .QN(n1530) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n3083), .CK(CLK), .QN(n1494) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n3082), .CK(CLK), .QN(n1458) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n3081), .CK(CLK), .QN(n1422) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n3080), .CK(CLK), .QN(n1386) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n3079), .CK(CLK), .QN(n1350) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n3078), .CK(CLK), .QN(n1314) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n3077), .CK(CLK), .QN(n1278) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n3076), .CK(CLK), .QN(n1242) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n3075), .CK(CLK), .QN(n1206) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n3074), .CK(CLK), .QN(n1170) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n3073), .CK(CLK), .QN(n1134) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n3072), .CK(CLK), .QN(n1098) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n3071), .CK(CLK), .QN(n1062) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n3070), .CK(CLK), .QN(n2194) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n3069), .CK(CLK), .QN(n2143) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n3068), .CK(CLK), .QN(n2107) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n3067), .CK(CLK), .QN(n2071) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n3066), .CK(CLK), .QN(n2035) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n3065), .CK(CLK), .QN(n1999) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n3064), .CK(CLK), .QN(n1963) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n3063), .CK(CLK), .QN(n1927) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n3062), .CK(CLK), .QN(n1891) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n3061), .CK(CLK), .QN(n1855) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n3060), .CK(CLK), .QN(n1819) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n3059), .CK(CLK), .QN(n1783) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n3058), .CK(CLK), .QN(n1747) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n3057), .CK(CLK), .QN(n1711) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n3056), .CK(CLK), .QN(n1675) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n3055), .CK(CLK), .QN(n1639) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n3054), .CK(CLK), .QN(n1603) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n3053), .CK(CLK), .QN(n1567) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n3052), .CK(CLK), .QN(n1531) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n3051), .CK(CLK), .QN(n1495) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n3050), .CK(CLK), .QN(n1459) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n3049), .CK(CLK), .QN(n1423) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n3048), .CK(CLK), .QN(n1387) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n3047), .CK(CLK), .QN(n1351) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n3046), .CK(CLK), .QN(n1315) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n3045), .CK(CLK), .QN(n1279) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n3044), .CK(CLK), .QN(n1243) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n3043), .CK(CLK), .QN(n1207) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n3042), .CK(CLK), .QN(n1171) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n3041), .CK(CLK), .QN(n1135) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n3040), .CK(CLK), .QN(n1099) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n3039), .CK(CLK), .QN(n1063) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n3038), .CK(CLK), .Q(n3773) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n3037), .CK(CLK), .Q(n3771) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n3036), .CK(CLK), .Q(n3770) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n3035), .CK(CLK), .Q(n3769) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n3034), .CK(CLK), .Q(n3768) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n3033), .CK(CLK), .Q(n3767) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n3032), .CK(CLK), .Q(n3766) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n3031), .CK(CLK), .Q(n3765) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n3030), .CK(CLK), .Q(n3764) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n3029), .CK(CLK), .Q(n3763) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n3028), .CK(CLK), .Q(n3762) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n3027), .CK(CLK), .Q(n3761) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n3026), .CK(CLK), .Q(n3760) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n3025), .CK(CLK), .Q(n3759) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n3024), .CK(CLK), .Q(n3758) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n3023), .CK(CLK), .Q(n3757) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n3022), .CK(CLK), .Q(n3756) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n3021), .CK(CLK), .Q(n3755) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n3020), .CK(CLK), .Q(n3754) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n3019), .CK(CLK), .Q(n3753) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n3018), .CK(CLK), .Q(n3752) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n3017), .CK(CLK), .Q(n3751) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n3016), .CK(CLK), .Q(n3750) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n3015), .CK(CLK), .Q(n3749) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n3014), .CK(CLK), .Q(n3748) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n3013), .CK(CLK), .Q(n3747) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n3012), .CK(CLK), .Q(n3746) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n3011), .CK(CLK), .Q(n3745) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n3010), .CK(CLK), .Q(n3744) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n3009), .CK(CLK), .Q(n3743) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n3008), .CK(CLK), .Q(n3742) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n3007), .CK(CLK), .Q(n3741) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n3006), .CK(CLK), .Q(n3739) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n3005), .CK(CLK), .Q(n3737) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n3004), .CK(CLK), .Q(n3736) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n3003), .CK(CLK), .Q(n3735) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n3002), .CK(CLK), .Q(n3734) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n3001), .CK(CLK), .Q(n3733) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n3000), .CK(CLK), .Q(n3732) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n2999), .CK(CLK), .Q(n3731) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n2998), .CK(CLK), .Q(n3730) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n2997), .CK(CLK), .Q(n3729) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n2996), .CK(CLK), .Q(n3728) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n2995), .CK(CLK), .Q(n3727) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n2994), .CK(CLK), .Q(n3726) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n2993), .CK(CLK), .Q(n3725) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n2992), .CK(CLK), .Q(n3724) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n2991), .CK(CLK), .Q(n3723) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n2990), .CK(CLK), .Q(n3722) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n2989), .CK(CLK), .Q(n3721) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n2988), .CK(CLK), .Q(n3720) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n2987), .CK(CLK), .Q(n3719) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n2986), .CK(CLK), .Q(n3718) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n2985), .CK(CLK), .Q(n3717) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n2984), .CK(CLK), .Q(n3716) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n2983), .CK(CLK), .Q(n3715) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n2982), .CK(CLK), .Q(n3714) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n2981), .CK(CLK), .Q(n3713) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n2980), .CK(CLK), .Q(n3712) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n2979), .CK(CLK), .Q(n3711) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n2978), .CK(CLK), .Q(n3710) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n2977), .CK(CLK), .Q(n3709) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n2976), .CK(CLK), .Q(n3708) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n2975), .CK(CLK), .Q(n3707) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n2974), .CK(CLK), .QN(n2187) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n2973), .CK(CLK), .QN(n2139) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n2972), .CK(CLK), .QN(n2103) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n2971), .CK(CLK), .QN(n2067) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n2970), .CK(CLK), .QN(n2031) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n2969), .CK(CLK), .QN(n1995) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n2968), .CK(CLK), .QN(n1959) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n2967), .CK(CLK), .QN(n1923) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n2966), .CK(CLK), .QN(n1887) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n2965), .CK(CLK), .QN(n1851) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n2964), .CK(CLK), .QN(n1815) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n2963), .CK(CLK), .QN(n1779) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n2962), .CK(CLK), .QN(n1743) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n2961), .CK(CLK), .QN(n1707) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n2960), .CK(CLK), .QN(n1671) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n2959), .CK(CLK), .QN(n1635) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n2958), .CK(CLK), .QN(n1599) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n2957), .CK(CLK), .QN(n1563) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n2956), .CK(CLK), .QN(n1527) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n2955), .CK(CLK), .QN(n1491) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n2954), .CK(CLK), .QN(n1455) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n2953), .CK(CLK), .QN(n1419) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n2952), .CK(CLK), .QN(n1383) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n2951), .CK(CLK), .QN(n1347) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n2950), .CK(CLK), .QN(n1311) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n2949), .CK(CLK), .QN(n1275) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n2948), .CK(CLK), .QN(n1239) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n2947), .CK(CLK), .QN(n1203) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n2946), .CK(CLK), .QN(n1167) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n2945), .CK(CLK), .QN(n1131) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n2944), .CK(CLK), .QN(n1095) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n2943), .CK(CLK), .QN(n1059) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n2942), .CK(CLK), .QN(n2189) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n2941), .CK(CLK), .QN(n2140) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n2940), .CK(CLK), .QN(n2104) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n2939), .CK(CLK), .QN(n2068) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n2938), .CK(CLK), .QN(n2032) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n2937), .CK(CLK), .QN(n1996) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n2936), .CK(CLK), .QN(n1960) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n2935), .CK(CLK), .QN(n1924) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n2934), .CK(CLK), .QN(n1888) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n2933), .CK(CLK), .QN(n1852) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n2932), .CK(CLK), .QN(n1816) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n2931), .CK(CLK), .QN(n1780) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n2930), .CK(CLK), .QN(n1744) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n2929), .CK(CLK), .QN(n1708) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n2928), .CK(CLK), .QN(n1672) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n2927), .CK(CLK), .QN(n1636) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n2926), .CK(CLK), .QN(n1600) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n2925), .CK(CLK), .QN(n1564) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n2924), .CK(CLK), .QN(n1528) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n2923), .CK(CLK), .QN(n1492) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n2922), .CK(CLK), .QN(n1456) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n2921), .CK(CLK), .QN(n1420) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n2920), .CK(CLK), .QN(n1384) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n2919), .CK(CLK), .QN(n1348) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n2918), .CK(CLK), .QN(n1312) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n2917), .CK(CLK), .QN(n1276) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n2916), .CK(CLK), .QN(n1240) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n2915), .CK(CLK), .QN(n1204) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n2914), .CK(CLK), .QN(n1168) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n2913), .CK(CLK), .QN(n1132) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n2912), .CK(CLK), .QN(n1096) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n2911), .CK(CLK), .QN(n1060) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n2910), .CK(CLK), .Q(n3637) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n2909), .CK(CLK), .Q(n3635) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n2908), .CK(CLK), .Q(n3634) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n2907), .CK(CLK), .Q(n3633) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n2906), .CK(CLK), .Q(n3632) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n2905), .CK(CLK), .Q(n3631) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n2904), .CK(CLK), .Q(n3630) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n2903), .CK(CLK), .Q(n3629) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n2902), .CK(CLK), .Q(n3628) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n2901), .CK(CLK), .Q(n3627) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n2900), .CK(CLK), .Q(n3626) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n2899), .CK(CLK), .Q(n3625) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n2898), .CK(CLK), .Q(n3624) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n2897), .CK(CLK), .Q(n3623) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n2896), .CK(CLK), .Q(n3622) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n2895), .CK(CLK), .Q(n3621) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n2894), .CK(CLK), .Q(n3620) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n2893), .CK(CLK), .Q(n3619) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n2892), .CK(CLK), .Q(n3618) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n2891), .CK(CLK), .Q(n3617) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n2890), .CK(CLK), .Q(n3616) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n2889), .CK(CLK), .Q(n3615) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n2888), .CK(CLK), .Q(n2526) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n2887), .CK(CLK), .Q(n2525) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n2886), .CK(CLK), .Q(n2524) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n2885), .CK(CLK), .Q(n2523) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n2884), .CK(CLK), .Q(n2522) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n2883), .CK(CLK), .Q(n2521) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n2882), .CK(CLK), .Q(n2520) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n2881), .CK(CLK), .Q(n2519) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n2880), .CK(CLK), .Q(n2518) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n2879), .CK(CLK), .Q(n2517) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n2878), .CK(CLK), .Q(n2515) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n2877), .CK(CLK), .Q(n2513) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n2876), .CK(CLK), .Q(n2512) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n2875), .CK(CLK), .Q(n2511) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n2874), .CK(CLK), .Q(n2510) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n2873), .CK(CLK), .Q(n2509) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n2872), .CK(CLK), .Q(n2508) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n2871), .CK(CLK), .Q(n2507) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n2870), .CK(CLK), .Q(n2506) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n2869), .CK(CLK), .Q(n2505) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n2868), .CK(CLK), .Q(n2504) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n2867), .CK(CLK), .Q(n2503) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n2866), .CK(CLK), .Q(n2502) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n2865), .CK(CLK), .Q(n2501) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n2864), .CK(CLK), .Q(n2500) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n2863), .CK(CLK), .Q(n2499) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n2862), .CK(CLK), .Q(n2498) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n2861), .CK(CLK), .Q(n2497) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n2860), .CK(CLK), .Q(n2496) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n2859), .CK(CLK), .Q(n2495) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n2858), .CK(CLK), .Q(n2494) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n2857), .CK(CLK), .Q(n2493) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n2856), .CK(CLK), .Q(n2492) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n2855), .CK(CLK), .Q(n2491) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n2854), .CK(CLK), .Q(n2490) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n2853), .CK(CLK), .Q(n2489) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n2852), .CK(CLK), .Q(n2488) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n2851), .CK(CLK), .Q(n2487) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n2850), .CK(CLK), .Q(n2486) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n2849), .CK(CLK), .Q(n2485) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n2848), .CK(CLK), .Q(n2484) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n2847), .CK(CLK), .Q(n2483) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n2846), .CK(CLK), .Q(n2481) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n2845), .CK(CLK), .Q(n2479) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n2844), .CK(CLK), .Q(n2478) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n2843), .CK(CLK), .Q(n2477) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n2842), .CK(CLK), .Q(n2476) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n2841), .CK(CLK), .Q(n2475) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n2840), .CK(CLK), .Q(n2474) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n2839), .CK(CLK), .Q(n2473) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n2838), .CK(CLK), .Q(n2472) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n2837), .CK(CLK), .Q(n2471) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n2836), .CK(CLK), .Q(n2470) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n2835), .CK(CLK), .Q(n2469) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n2834), .CK(CLK), .Q(n2468) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n2833), .CK(CLK), .Q(n2467) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n2832), .CK(CLK), .Q(n2466) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n2831), .CK(CLK), .Q(n2465) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n2830), .CK(CLK), .Q(n2464) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n2829), .CK(CLK), .Q(n2463) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n2828), .CK(CLK), .Q(n2462) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n2827), .CK(CLK), .Q(n2461) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n2826), .CK(CLK), .Q(n2460) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n2825), .CK(CLK), .Q(n2459) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n2824), .CK(CLK), .Q(n2458) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n2823), .CK(CLK), .Q(n2457) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n2822), .CK(CLK), .Q(n2456) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n2821), .CK(CLK), .Q(n2455) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n2820), .CK(CLK), .Q(n2454) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n2819), .CK(CLK), .Q(n2453) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n2818), .CK(CLK), .Q(n2452) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n2817), .CK(CLK), .Q(n2451) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n2816), .CK(CLK), .Q(n2450) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n2815), .CK(CLK), .Q(n2449) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n2814), .CK(CLK), .Q(n2443) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n2813), .CK(CLK), .Q(n2441) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n2812), .CK(CLK), .Q(n2440) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n2811), .CK(CLK), .Q(n2439) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n2810), .CK(CLK), .Q(n2438) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n2809), .CK(CLK), .Q(n2437) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n2808), .CK(CLK), .Q(n2436) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n2807), .CK(CLK), .Q(n2435) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n2806), .CK(CLK), .Q(n2434) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n2805), .CK(CLK), .Q(n2433) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n2804), .CK(CLK), .Q(n2432) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n2803), .CK(CLK), .Q(n2431) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n2802), .CK(CLK), .Q(n2430) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n2801), .CK(CLK), .Q(n2429) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n2800), .CK(CLK), .Q(n2428) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n2799), .CK(CLK), .Q(n2427) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n2798), .CK(CLK), .Q(n2426) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n2797), .CK(CLK), .Q(n2425) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n2796), .CK(CLK), .Q(n2424) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n2795), .CK(CLK), .Q(n2423) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n2794), .CK(CLK), .Q(n2422) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n2793), .CK(CLK), .Q(n2421) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n2792), .CK(CLK), .Q(n2420) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n2791), .CK(CLK), .Q(n2419) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n2790), .CK(CLK), .Q(n2418) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n2789), .CK(CLK), .Q(n2417) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n2788), .CK(CLK), .Q(n2416) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n2787), .CK(CLK), .Q(n2415) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n2786), .CK(CLK), .Q(n2414) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n2785), .CK(CLK), .Q(n2413) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n2784), .CK(CLK), .Q(n2412) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n2783), .CK(CLK), .Q(n2411) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n2782), .CK(CLK), .QN(n2182) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n2781), .CK(CLK), .QN(n2136) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n2780), .CK(CLK), .QN(n2100) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n2779), .CK(CLK), .QN(n2064) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n2778), .CK(CLK), .QN(n2028) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n2777), .CK(CLK), .QN(n1992) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n2776), .CK(CLK), .QN(n1956) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n2775), .CK(CLK), .QN(n1920) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n2774), .CK(CLK), .QN(n1884) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n2773), .CK(CLK), .QN(n1848) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n2772), .CK(CLK), .QN(n1812) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n2771), .CK(CLK), .QN(n1776) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n2770), .CK(CLK), .QN(n1740) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n2769), .CK(CLK), .QN(n1704) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n2768), .CK(CLK), .QN(n1668) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n2767), .CK(CLK), .QN(n1632) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n2766), .CK(CLK), .QN(n1596) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n2765), .CK(CLK), .QN(n1560) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n2764), .CK(CLK), .QN(n1524) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n2763), .CK(CLK), .QN(n1488) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n2762), .CK(CLK), .QN(n1452) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n2761), .CK(CLK), .QN(n1416) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n2760), .CK(CLK), .QN(n1380) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n2759), .CK(CLK), .QN(n1344) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n2758), .CK(CLK), .QN(n1308) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n2757), .CK(CLK), .QN(n1272) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n2756), .CK(CLK), .QN(n1236) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n2755), .CK(CLK), .QN(n1200) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n2754), .CK(CLK), .QN(n1164) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n2753), .CK(CLK), .QN(n1128) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n2752), .CK(CLK), .QN(n1092) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n2751), .CK(CLK), .QN(n1054) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n2750), .CK(CLK), .QN(n2184) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n2749), .CK(CLK), .QN(n2137) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n2748), .CK(CLK), .QN(n2101) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n2747), .CK(CLK), .QN(n2065) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n2746), .CK(CLK), .QN(n2029) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n2745), .CK(CLK), .QN(n1993) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n2744), .CK(CLK), .QN(n1957) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n2743), .CK(CLK), .QN(n1921) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n2742), .CK(CLK), .QN(n1885) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n2741), .CK(CLK), .QN(n1849) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n2740), .CK(CLK), .QN(n1813) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n2739), .CK(CLK), .QN(n1777) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n2738), .CK(CLK), .QN(n1741) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n2737), .CK(CLK), .QN(n1705) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n2736), .CK(CLK), .QN(n1669) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n2735), .CK(CLK), .QN(n1633) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n2734), .CK(CLK), .QN(n1597) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n2733), .CK(CLK), .QN(n1561) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n2732), .CK(CLK), .QN(n1525) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n2731), .CK(CLK), .QN(n1489) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n2730), .CK(CLK), .QN(n1453) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n2729), .CK(CLK), .QN(n1417) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n2728), .CK(CLK), .QN(n1381) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n2727), .CK(CLK), .QN(n1345) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n2726), .CK(CLK), .QN(n1309) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n2725), .CK(CLK), .QN(n1273) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n2724), .CK(CLK), .QN(n1237) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n2723), .CK(CLK), .QN(n1201) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n2722), .CK(CLK), .QN(n1165) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n2721), .CK(CLK), .QN(n1129) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n2720), .CK(CLK), .QN(n1093) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n2719), .CK(CLK), .QN(n1055) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n2718), .CK(CLK), .Q(n2341) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n2717), .CK(CLK), .Q(n2339) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n2716), .CK(CLK), .Q(n2338) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n2715), .CK(CLK), .Q(n2337) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n2714), .CK(CLK), .Q(n2336) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n2713), .CK(CLK), .Q(n2335) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n2712), .CK(CLK), .Q(n2334) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n2711), .CK(CLK), .Q(n2333) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n2710), .CK(CLK), .Q(n2332) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n2709), .CK(CLK), .Q(n2331) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n2708), .CK(CLK), .Q(n2330) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n2707), .CK(CLK), .Q(n2329) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n2706), .CK(CLK), .Q(n2328) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n2705), .CK(CLK), .Q(n2327) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n2704), .CK(CLK), .Q(n2326) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n2703), .CK(CLK), .Q(n2325) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n2702), .CK(CLK), .Q(n2324) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n2701), .CK(CLK), .Q(n2323) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n2700), .CK(CLK), .Q(n2322) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n2699), .CK(CLK), .Q(n2321) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n2698), .CK(CLK), .Q(n2320) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n2697), .CK(CLK), .Q(n2319) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n2696), .CK(CLK), .Q(n2318) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n2695), .CK(CLK), .Q(n2317) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n2694), .CK(CLK), .Q(n2316) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n2693), .CK(CLK), .Q(n2315) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n2692), .CK(CLK), .Q(n2314) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n2691), .CK(CLK), .Q(n2313) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n2690), .CK(CLK), .Q(n2312) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n2689), .CK(CLK), .Q(n2311) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n2688), .CK(CLK), .Q(n2310) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n2687), .CK(CLK), .Q(n2309) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n2686), .CK(CLK), .Q(n2307) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n2685), .CK(CLK), .Q(n2305) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n2684), .CK(CLK), .Q(n2304) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n2683), .CK(CLK), .Q(n2303) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n2682), .CK(CLK), .Q(n2302) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n2681), .CK(CLK), .Q(n2301) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n2680), .CK(CLK), .Q(n2300) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n2679), .CK(CLK), .Q(n2299) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n2678), .CK(CLK), .Q(n2298) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n2677), .CK(CLK), .Q(n2297) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n2676), .CK(CLK), .Q(n2296) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n2675), .CK(CLK), .Q(n2295) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n2674), .CK(CLK), .Q(n2294) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n2673), .CK(CLK), .Q(n2293) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n2672), .CK(CLK), .Q(n2292) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n2671), .CK(CLK), .Q(n2291) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n2670), .CK(CLK), .Q(n2290) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n2669), .CK(CLK), .Q(n2289) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n2668), .CK(CLK), .Q(n2288) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n2667), .CK(CLK), .Q(n2287) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n2666), .CK(CLK), .Q(n2286) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n2665), .CK(CLK), .Q(n2285) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n2664), .CK(CLK), .Q(n2284) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n2663), .CK(CLK), .Q(n2283) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n2662), .CK(CLK), .Q(n2282) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n2661), .CK(CLK), .Q(n2281) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n2660), .CK(CLK), .Q(n2280) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n2659), .CK(CLK), .Q(n2279) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n2658), .CK(CLK), .Q(n2278) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n2657), .CK(CLK), .Q(n2277) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n2656), .CK(CLK), .Q(n2276) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n2655), .CK(CLK), .Q(n2275) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n2654), .CK(CLK), .QN(n2177) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n2653), .CK(CLK), .QN(n2133) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n2652), .CK(CLK), .QN(n2097) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n2651), .CK(CLK), .QN(n2061) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n2650), .CK(CLK), .QN(n2025) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n2649), .CK(CLK), .QN(n1989) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n2648), .CK(CLK), .QN(n1953) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n2647), .CK(CLK), .QN(n1917) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n2646), .CK(CLK), .QN(n1881) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n2645), .CK(CLK), .QN(n1845) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n2644), .CK(CLK), .QN(n1809) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n2643), .CK(CLK), .QN(n1773) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n2642), .CK(CLK), .QN(n1737) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n2641), .CK(CLK), .QN(n1701) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n2640), .CK(CLK), .QN(n1665) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n2639), .CK(CLK), .QN(n1629) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n2638), .CK(CLK), .QN(n1593) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n2637), .CK(CLK), .QN(n1557) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n2636), .CK(CLK), .QN(n1521) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n2635), .CK(CLK), .QN(n1485) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n2634), .CK(CLK), .QN(n1449) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n2633), .CK(CLK), .QN(n1413) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n2632), .CK(CLK), .QN(n1377) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n2631), .CK(CLK), .QN(n1341) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n2630), .CK(CLK), .QN(n1305) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n2629), .CK(CLK), .QN(n1269) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n2628), .CK(CLK), .QN(n1233) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n2627), .CK(CLK), .QN(n1197) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n2626), .CK(CLK), .QN(n1161) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n2625), .CK(CLK), .QN(n1125) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n2624), .CK(CLK), .QN(n1089) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n2623), .CK(CLK), .QN(n1051) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n2622), .CK(CLK), .QN(n2179) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n2621), .CK(CLK), .QN(n2134) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n2620), .CK(CLK), .QN(n2098) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n2619), .CK(CLK), .QN(n2062) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n2618), .CK(CLK), .QN(n2026) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n2617), .CK(CLK), .QN(n1990) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n2616), .CK(CLK), .QN(n1954) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n2615), .CK(CLK), .QN(n1918) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n2614), .CK(CLK), .QN(n1882) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n2613), .CK(CLK), .QN(n1846) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n2612), .CK(CLK), .QN(n1810) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n2611), .CK(CLK), .QN(n1774) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n2610), .CK(CLK), .QN(n1738) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n2609), .CK(CLK), .QN(n1702) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n2608), .CK(CLK), .QN(n1666) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n2607), .CK(CLK), .QN(n1630) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n2606), .CK(CLK), .QN(n1594) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n2605), .CK(CLK), .QN(n1558) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n2604), .CK(CLK), .QN(n1522) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n2603), .CK(CLK), .QN(n1486) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n2602), .CK(CLK), .QN(n1450) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n2601), .CK(CLK), .QN(n1414) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n2600), .CK(CLK), .QN(n1378) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n2599), .CK(CLK), .QN(n1342) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n2598), .CK(CLK), .QN(n1306) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n2597), .CK(CLK), .QN(n1270) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n2596), .CK(CLK), .QN(n1234) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n2595), .CK(CLK), .QN(n1198) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n2594), .CK(CLK), .QN(n1162) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n2593), .CK(CLK), .QN(n1126) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n2592), .CK(CLK), .QN(n1090) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n2591), .CK(CLK), .QN(n1052) );
  DFF_X1 \OUT1_reg[13]  ( .D(n2572), .CK(CLK), .Q(OUT1[13]), .QN(n1540) );
  DFF_X1 \OUT1_reg[12]  ( .D(n2571), .CK(CLK), .Q(OUT1[12]), .QN(n1504) );
  DFF_X1 \OUT1_reg[11]  ( .D(n2570), .CK(CLK), .Q(OUT1[11]), .QN(n1468) );
  DFF_X1 \OUT2_reg[23]  ( .D(n2550), .CK(CLK), .Q(OUT2[23]), .QN(n854) );
  DFF_X1 \OUT2_reg[22]  ( .D(n2549), .CK(CLK), .Q(OUT2[22]), .QN(n834) );
  DFF_X1 \OUT2_reg[21]  ( .D(n2548), .CK(CLK), .Q(OUT2[21]), .QN(n814) );
  DFF_X1 \OUT2_reg[20]  ( .D(n2547), .CK(CLK), .Q(OUT2[20]), .QN(n794) );
  DFF_X1 \OUT2_reg[19]  ( .D(n2546), .CK(CLK), .Q(OUT2[19]), .QN(n774) );
  DFF_X1 \OUT2_reg[18]  ( .D(n2545), .CK(CLK), .Q(OUT2[18]), .QN(n754) );
  DFF_X1 \OUT2_reg[17]  ( .D(n2544), .CK(CLK), .Q(OUT2[17]), .QN(n734) );
  DFF_X1 \OUT2_reg[16]  ( .D(n2543), .CK(CLK), .Q(OUT2[16]), .QN(n714) );
  DFF_X1 \OUT2_reg[15]  ( .D(n2542), .CK(CLK), .Q(OUT2[15]), .QN(n694) );
  DFF_X1 \OUT2_reg[14]  ( .D(n2541), .CK(CLK), .Q(OUT2[14]), .QN(n674) );
  DFF_X1 \OUT2_reg[13]  ( .D(n2540), .CK(CLK), .Q(OUT2[13]), .QN(n654) );
  DFF_X1 \OUT2_reg[12]  ( .D(n2539), .CK(CLK), .Q(OUT2[12]), .QN(n634) );
  DFF_X1 \OUT2_reg[11]  ( .D(n2538), .CK(CLK), .Q(OUT2[11]), .QN(n614) );
  DFF_X1 \OUT2_reg[10]  ( .D(n2537), .CK(CLK), .Q(OUT2[10]), .QN(n594) );
  DFF_X1 \OUT2_reg[9]  ( .D(n2536), .CK(CLK), .Q(OUT2[9]), .QN(n574) );
  DFF_X1 \OUT2_reg[8]  ( .D(n2535), .CK(CLK), .Q(OUT2[8]), .QN(n554) );
  DFF_X1 \OUT2_reg[7]  ( .D(n2534), .CK(CLK), .Q(OUT2[7]), .QN(n534) );
  DFF_X1 \OUT2_reg[6]  ( .D(n2533), .CK(CLK), .Q(OUT2[6]), .QN(n514) );
  DFF_X1 \OUT2_reg[5]  ( .D(n2532), .CK(CLK), .Q(OUT2[5]), .QN(n494) );
  DFF_X1 \OUT2_reg[4]  ( .D(n2531), .CK(CLK), .Q(OUT2[4]), .QN(n474) );
  DFF_X1 \OUT2_reg[3]  ( .D(n2530), .CK(CLK), .Q(OUT2[3]), .QN(n454) );
  DFF_X1 \OUT2_reg[2]  ( .D(n2529), .CK(CLK), .Q(OUT2[2]), .QN(n434) );
  DFF_X1 \OUT2_reg[1]  ( .D(n2528), .CK(CLK), .Q(OUT2[1]), .QN(n414) );
  DFF_X1 \OUT2_reg[0]  ( .D(n2527), .CK(CLK), .Q(OUT2[0]), .QN(n394) );
  AND2_X1 U3 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n1) );
  AND2_X1 U4 ( .A1(ADD_RD2[1]), .A2(n371), .ZN(n2) );
  AND2_X1 U5 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n3) );
  AND2_X1 U6 ( .A1(ADD_RD1[1]), .A2(n1035), .ZN(n4) );
  CLKBUF_X3 U7 ( .A(n1031), .Z(n162) );
  CLKBUF_X3 U8 ( .A(n2205), .Z(n264) );
  BUF_X1 U9 ( .A(n3806), .Z(n309) );
  BUF_X1 U10 ( .A(n3806), .Z(n310) );
  BUF_X1 U11 ( .A(n2374), .Z(n279) );
  BUF_X1 U12 ( .A(n2374), .Z(n280) );
  BUF_X1 U13 ( .A(n2408), .Z(n282) );
  BUF_X1 U14 ( .A(n2408), .Z(n283) );
  BUF_X1 U15 ( .A(n3670), .Z(n297) );
  BUF_X1 U16 ( .A(n3670), .Z(n298) );
  BUF_X1 U17 ( .A(n3704), .Z(n300) );
  BUF_X1 U18 ( .A(n3704), .Z(n301) );
  BUF_X1 U19 ( .A(n3841), .Z(n312) );
  BUF_X1 U20 ( .A(n3841), .Z(n313) );
  BUF_X1 U21 ( .A(n2238), .Z(n267) );
  BUF_X1 U22 ( .A(n2238), .Z(n268) );
  BUF_X1 U23 ( .A(n2272), .Z(n270) );
  BUF_X1 U24 ( .A(n2272), .Z(n271) );
  BUF_X1 U25 ( .A(n2442), .Z(n285) );
  BUF_X1 U26 ( .A(n2442), .Z(n286) );
  BUF_X1 U27 ( .A(n2306), .Z(n273) );
  BUF_X1 U28 ( .A(n2306), .Z(n274) );
  BUF_X1 U29 ( .A(n2340), .Z(n276) );
  BUF_X1 U30 ( .A(n2340), .Z(n277) );
  BUF_X1 U31 ( .A(n2480), .Z(n288) );
  BUF_X1 U32 ( .A(n2480), .Z(n289) );
  BUF_X1 U33 ( .A(n3738), .Z(n303) );
  BUF_X1 U34 ( .A(n3738), .Z(n304) );
  BUF_X1 U35 ( .A(n3772), .Z(n306) );
  BUF_X1 U36 ( .A(n3772), .Z(n307) );
  BUF_X1 U37 ( .A(n2514), .Z(n291) );
  BUF_X1 U38 ( .A(n2514), .Z(n292) );
  BUF_X1 U39 ( .A(n3636), .Z(n294) );
  BUF_X1 U40 ( .A(n3636), .Z(n295) );
  BUF_X1 U41 ( .A(n7), .Z(n159) );
  BUF_X1 U42 ( .A(n7), .Z(n160) );
  BUF_X1 U43 ( .A(n8), .Z(n261) );
  BUF_X1 U44 ( .A(n8), .Z(n262) );
  BUF_X1 U45 ( .A(n2169), .Z(n201) );
  BUF_X1 U46 ( .A(n2169), .Z(n202) );
  BUF_X1 U47 ( .A(n5), .Z(n129) );
  BUF_X1 U48 ( .A(n5), .Z(n130) );
  BUF_X1 U49 ( .A(n6), .Z(n231) );
  BUF_X1 U50 ( .A(n6), .Z(n232) );
  BUF_X1 U51 ( .A(n1004), .Z(n99) );
  BUF_X1 U52 ( .A(n1004), .Z(n100) );
  BUF_X1 U53 ( .A(n3806), .Z(n311) );
  BUF_X1 U54 ( .A(n2374), .Z(n281) );
  BUF_X1 U55 ( .A(n2408), .Z(n284) );
  BUF_X1 U56 ( .A(n3670), .Z(n299) );
  BUF_X1 U57 ( .A(n3704), .Z(n302) );
  BUF_X1 U58 ( .A(n3841), .Z(n314) );
  BUF_X1 U59 ( .A(n2238), .Z(n269) );
  BUF_X1 U60 ( .A(n2272), .Z(n272) );
  BUF_X1 U61 ( .A(n2442), .Z(n287) );
  BUF_X1 U62 ( .A(n2306), .Z(n275) );
  BUF_X1 U63 ( .A(n2340), .Z(n278) );
  BUF_X1 U64 ( .A(n2480), .Z(n290) );
  BUF_X1 U65 ( .A(n3738), .Z(n305) );
  BUF_X1 U66 ( .A(n3772), .Z(n308) );
  BUF_X1 U67 ( .A(n2514), .Z(n293) );
  BUF_X1 U68 ( .A(n3636), .Z(n296) );
  BUF_X1 U69 ( .A(n7), .Z(n161) );
  BUF_X1 U70 ( .A(n8), .Z(n263) );
  BUF_X1 U71 ( .A(n2169), .Z(n203) );
  BUF_X1 U72 ( .A(n5), .Z(n131) );
  BUF_X1 U73 ( .A(n6), .Z(n233) );
  BUF_X1 U74 ( .A(n1004), .Z(n101) );
  BUF_X1 U75 ( .A(n4221), .Z(n345) );
  BUF_X1 U76 ( .A(n4221), .Z(n346) );
  BUF_X1 U77 ( .A(n4256), .Z(n348) );
  BUF_X1 U78 ( .A(n4256), .Z(n349) );
  BUF_X1 U79 ( .A(n4393), .Z(n357) );
  BUF_X1 U80 ( .A(n4393), .Z(n358) );
  BUF_X1 U81 ( .A(n4460), .Z(n360) );
  BUF_X1 U82 ( .A(n4460), .Z(n361) );
  BUF_X1 U83 ( .A(n3943), .Z(n321) );
  BUF_X1 U84 ( .A(n3943), .Z(n322) );
  BUF_X1 U85 ( .A(n3977), .Z(n324) );
  BUF_X1 U86 ( .A(n3977), .Z(n325) );
  BUF_X1 U87 ( .A(n4079), .Z(n333) );
  BUF_X1 U88 ( .A(n4079), .Z(n334) );
  BUF_X1 U89 ( .A(n4114), .Z(n336) );
  BUF_X1 U90 ( .A(n4114), .Z(n337) );
  BUF_X1 U91 ( .A(n4151), .Z(n339) );
  BUF_X1 U92 ( .A(n4151), .Z(n340) );
  BUF_X1 U93 ( .A(n4186), .Z(n342) );
  BUF_X1 U94 ( .A(n4186), .Z(n343) );
  BUF_X1 U95 ( .A(n4291), .Z(n351) );
  BUF_X1 U96 ( .A(n4291), .Z(n352) );
  BUF_X1 U97 ( .A(n4357), .Z(n354) );
  BUF_X1 U98 ( .A(n4357), .Z(n355) );
  BUF_X1 U99 ( .A(n3875), .Z(n315) );
  BUF_X1 U100 ( .A(n3875), .Z(n316) );
  BUF_X1 U101 ( .A(n3909), .Z(n318) );
  BUF_X1 U102 ( .A(n3909), .Z(n319) );
  BUF_X1 U103 ( .A(n4011), .Z(n327) );
  BUF_X1 U104 ( .A(n4011), .Z(n328) );
  BUF_X1 U105 ( .A(n4045), .Z(n330) );
  BUF_X1 U106 ( .A(n4045), .Z(n331) );
  BUF_X1 U107 ( .A(n2190), .Z(n240) );
  BUF_X1 U108 ( .A(n2190), .Z(n241) );
  BUF_X1 U109 ( .A(n2195), .Z(n252) );
  BUF_X1 U110 ( .A(n2195), .Z(n253) );
  BUF_X1 U111 ( .A(n2161), .Z(n180) );
  BUF_X1 U112 ( .A(n2161), .Z(n181) );
  BUF_X1 U113 ( .A(n2166), .Z(n192) );
  BUF_X1 U114 ( .A(n2166), .Z(n193) );
  BUF_X1 U115 ( .A(n2171), .Z(n204) );
  BUF_X1 U116 ( .A(n2171), .Z(n205) );
  BUF_X1 U117 ( .A(n2156), .Z(n168) );
  BUF_X1 U118 ( .A(n2156), .Z(n169) );
  BUF_X1 U119 ( .A(n2185), .Z(n228) );
  BUF_X1 U120 ( .A(n2185), .Z(n229) );
  BUF_X1 U121 ( .A(n2180), .Z(n216) );
  BUF_X1 U122 ( .A(n2180), .Z(n217) );
  BUF_X1 U123 ( .A(n2188), .Z(n237) );
  BUF_X1 U124 ( .A(n2188), .Z(n238) );
  BUF_X1 U125 ( .A(n2193), .Z(n249) );
  BUF_X1 U126 ( .A(n2193), .Z(n250) );
  BUF_X1 U127 ( .A(n2159), .Z(n177) );
  BUF_X1 U128 ( .A(n2159), .Z(n178) );
  BUF_X1 U129 ( .A(n2164), .Z(n189) );
  BUF_X1 U130 ( .A(n2164), .Z(n190) );
  BUF_X1 U131 ( .A(n2154), .Z(n165) );
  BUF_X1 U132 ( .A(n2154), .Z(n166) );
  BUF_X1 U133 ( .A(n2183), .Z(n225) );
  BUF_X1 U134 ( .A(n2183), .Z(n226) );
  BUF_X1 U135 ( .A(n2178), .Z(n213) );
  BUF_X1 U136 ( .A(n2178), .Z(n214) );
  BUF_X1 U137 ( .A(n27), .Z(n141) );
  BUF_X1 U138 ( .A(n27), .Z(n142) );
  BUF_X1 U139 ( .A(n28), .Z(n153) );
  BUF_X1 U140 ( .A(n28), .Z(n154) );
  BUF_X1 U141 ( .A(n29), .Z(n81) );
  BUF_X1 U142 ( .A(n29), .Z(n82) );
  BUF_X1 U143 ( .A(n30), .Z(n93) );
  BUF_X1 U144 ( .A(n30), .Z(n94) );
  BUF_X1 U145 ( .A(n31), .Z(n105) );
  BUF_X1 U146 ( .A(n31), .Z(n106) );
  BUF_X1 U147 ( .A(n19), .Z(n117) );
  BUF_X1 U148 ( .A(n19), .Z(n118) );
  BUF_X1 U149 ( .A(n32), .Z(n243) );
  BUF_X1 U150 ( .A(n32), .Z(n244) );
  BUF_X1 U151 ( .A(n33), .Z(n69) );
  BUF_X1 U152 ( .A(n33), .Z(n70) );
  BUF_X1 U153 ( .A(n34), .Z(n255) );
  BUF_X1 U154 ( .A(n34), .Z(n256) );
  BUF_X1 U155 ( .A(n35), .Z(n183) );
  BUF_X1 U156 ( .A(n35), .Z(n184) );
  BUF_X1 U157 ( .A(n36), .Z(n195) );
  BUF_X1 U158 ( .A(n36), .Z(n196) );
  BUF_X1 U159 ( .A(n37), .Z(n207) );
  BUF_X1 U160 ( .A(n37), .Z(n208) );
  BUF_X1 U161 ( .A(n20), .Z(n219) );
  BUF_X1 U162 ( .A(n20), .Z(n220) );
  BUF_X1 U163 ( .A(n38), .Z(n171) );
  BUF_X1 U164 ( .A(n38), .Z(n172) );
  BUF_X1 U165 ( .A(n1017), .Z(n135) );
  BUF_X1 U166 ( .A(n1017), .Z(n136) );
  BUF_X1 U167 ( .A(n1020), .Z(n147) );
  BUF_X1 U168 ( .A(n1020), .Z(n148) );
  BUF_X1 U169 ( .A(n998), .Z(n75) );
  BUF_X1 U170 ( .A(n998), .Z(n76) );
  BUF_X1 U171 ( .A(n1001), .Z(n87) );
  BUF_X1 U172 ( .A(n1001), .Z(n88) );
  BUF_X1 U173 ( .A(n995), .Z(n63) );
  BUF_X1 U174 ( .A(n995), .Z(n64) );
  BUF_X1 U175 ( .A(n1014), .Z(n123) );
  BUF_X1 U176 ( .A(n1014), .Z(n124) );
  BUF_X1 U177 ( .A(n1011), .Z(n111) );
  BUF_X1 U178 ( .A(n1011), .Z(n112) );
  BUF_X1 U179 ( .A(n1018), .Z(n138) );
  BUF_X1 U180 ( .A(n1018), .Z(n139) );
  BUF_X1 U181 ( .A(n1021), .Z(n150) );
  BUF_X1 U182 ( .A(n1021), .Z(n151) );
  BUF_X1 U183 ( .A(n999), .Z(n78) );
  BUF_X1 U184 ( .A(n999), .Z(n79) );
  BUF_X1 U185 ( .A(n1002), .Z(n90) );
  BUF_X1 U186 ( .A(n1002), .Z(n91) );
  BUF_X1 U187 ( .A(n1005), .Z(n102) );
  BUF_X1 U188 ( .A(n1005), .Z(n103) );
  BUF_X1 U189 ( .A(n996), .Z(n66) );
  BUF_X1 U190 ( .A(n996), .Z(n67) );
  BUF_X1 U191 ( .A(n1015), .Z(n126) );
  BUF_X1 U192 ( .A(n1015), .Z(n127) );
  BUF_X1 U193 ( .A(n1012), .Z(n114) );
  BUF_X1 U194 ( .A(n1012), .Z(n115) );
  BUF_X1 U195 ( .A(n21), .Z(n144) );
  BUF_X1 U196 ( .A(n21), .Z(n145) );
  BUF_X1 U197 ( .A(n22), .Z(n156) );
  BUF_X1 U198 ( .A(n22), .Z(n157) );
  BUF_X1 U199 ( .A(n17), .Z(n132) );
  BUF_X1 U200 ( .A(n17), .Z(n133) );
  BUF_X1 U201 ( .A(n42), .Z(n84) );
  BUF_X1 U202 ( .A(n42), .Z(n85) );
  BUF_X1 U203 ( .A(n40), .Z(n96) );
  BUF_X1 U204 ( .A(n40), .Z(n97) );
  BUF_X1 U205 ( .A(n43), .Z(n108) );
  BUF_X1 U206 ( .A(n43), .Z(n109) );
  BUF_X1 U207 ( .A(n15), .Z(n120) );
  BUF_X1 U208 ( .A(n15), .Z(n121) );
  BUF_X1 U209 ( .A(n23), .Z(n72) );
  BUF_X1 U210 ( .A(n23), .Z(n73) );
  BUF_X1 U211 ( .A(n24), .Z(n246) );
  BUF_X1 U212 ( .A(n24), .Z(n247) );
  BUF_X1 U213 ( .A(n18), .Z(n234) );
  BUF_X1 U214 ( .A(n18), .Z(n235) );
  BUF_X1 U215 ( .A(n25), .Z(n258) );
  BUF_X1 U216 ( .A(n25), .Z(n259) );
  BUF_X1 U217 ( .A(n44), .Z(n186) );
  BUF_X1 U218 ( .A(n44), .Z(n187) );
  BUF_X1 U219 ( .A(n41), .Z(n198) );
  BUF_X1 U220 ( .A(n41), .Z(n199) );
  BUF_X1 U221 ( .A(n16), .Z(n222) );
  BUF_X1 U222 ( .A(n16), .Z(n223) );
  BUF_X1 U223 ( .A(n45), .Z(n210) );
  BUF_X1 U224 ( .A(n45), .Z(n211) );
  BUF_X1 U225 ( .A(n26), .Z(n174) );
  BUF_X1 U226 ( .A(n26), .Z(n175) );
  BUF_X1 U227 ( .A(n4221), .Z(n347) );
  BUF_X1 U228 ( .A(n4256), .Z(n350) );
  BUF_X1 U229 ( .A(n4393), .Z(n359) );
  BUF_X1 U230 ( .A(n4460), .Z(n362) );
  BUF_X1 U231 ( .A(n3943), .Z(n323) );
  BUF_X1 U232 ( .A(n3977), .Z(n326) );
  BUF_X1 U233 ( .A(n4079), .Z(n335) );
  BUF_X1 U234 ( .A(n4114), .Z(n338) );
  BUF_X1 U235 ( .A(n4151), .Z(n341) );
  BUF_X1 U236 ( .A(n4186), .Z(n344) );
  BUF_X1 U237 ( .A(n4291), .Z(n353) );
  BUF_X1 U238 ( .A(n4357), .Z(n356) );
  BUF_X1 U239 ( .A(n3875), .Z(n317) );
  BUF_X1 U240 ( .A(n3909), .Z(n320) );
  BUF_X1 U241 ( .A(n4045), .Z(n332) );
  BUF_X1 U242 ( .A(n4011), .Z(n329) );
  BUF_X1 U243 ( .A(n2190), .Z(n242) );
  BUF_X1 U244 ( .A(n2195), .Z(n254) );
  BUF_X1 U245 ( .A(n2161), .Z(n182) );
  BUF_X1 U246 ( .A(n2166), .Z(n194) );
  BUF_X1 U247 ( .A(n2171), .Z(n206) );
  BUF_X1 U248 ( .A(n2156), .Z(n170) );
  BUF_X1 U249 ( .A(n2185), .Z(n230) );
  BUF_X1 U250 ( .A(n2180), .Z(n218) );
  BUF_X1 U251 ( .A(n2188), .Z(n239) );
  BUF_X1 U252 ( .A(n2193), .Z(n251) );
  BUF_X1 U253 ( .A(n2159), .Z(n179) );
  BUF_X1 U254 ( .A(n2164), .Z(n191) );
  BUF_X1 U255 ( .A(n2154), .Z(n167) );
  BUF_X1 U256 ( .A(n2183), .Z(n227) );
  BUF_X1 U257 ( .A(n2178), .Z(n215) );
  BUF_X1 U258 ( .A(n27), .Z(n143) );
  BUF_X1 U259 ( .A(n28), .Z(n155) );
  BUF_X1 U260 ( .A(n29), .Z(n83) );
  BUF_X1 U261 ( .A(n30), .Z(n95) );
  BUF_X1 U262 ( .A(n31), .Z(n107) );
  BUF_X1 U263 ( .A(n19), .Z(n119) );
  BUF_X1 U264 ( .A(n32), .Z(n245) );
  BUF_X1 U265 ( .A(n33), .Z(n71) );
  BUF_X1 U266 ( .A(n34), .Z(n257) );
  BUF_X1 U267 ( .A(n35), .Z(n185) );
  BUF_X1 U268 ( .A(n36), .Z(n197) );
  BUF_X1 U269 ( .A(n37), .Z(n209) );
  BUF_X1 U270 ( .A(n20), .Z(n221) );
  BUF_X1 U271 ( .A(n38), .Z(n173) );
  BUF_X1 U272 ( .A(n1017), .Z(n137) );
  BUF_X1 U273 ( .A(n1020), .Z(n149) );
  BUF_X1 U274 ( .A(n998), .Z(n77) );
  BUF_X1 U275 ( .A(n1001), .Z(n89) );
  BUF_X1 U276 ( .A(n995), .Z(n65) );
  BUF_X1 U277 ( .A(n1014), .Z(n125) );
  BUF_X1 U278 ( .A(n1011), .Z(n113) );
  BUF_X1 U279 ( .A(n1018), .Z(n140) );
  BUF_X1 U280 ( .A(n1021), .Z(n152) );
  BUF_X1 U281 ( .A(n999), .Z(n80) );
  BUF_X1 U282 ( .A(n1002), .Z(n92) );
  BUF_X1 U283 ( .A(n1005), .Z(n104) );
  BUF_X1 U284 ( .A(n996), .Z(n68) );
  BUF_X1 U285 ( .A(n1015), .Z(n128) );
  BUF_X1 U286 ( .A(n1012), .Z(n116) );
  BUF_X1 U287 ( .A(n21), .Z(n146) );
  BUF_X1 U288 ( .A(n22), .Z(n158) );
  BUF_X1 U289 ( .A(n17), .Z(n134) );
  BUF_X1 U290 ( .A(n42), .Z(n86) );
  BUF_X1 U291 ( .A(n40), .Z(n98) );
  BUF_X1 U292 ( .A(n43), .Z(n110) );
  BUF_X1 U293 ( .A(n15), .Z(n122) );
  BUF_X1 U294 ( .A(n23), .Z(n74) );
  BUF_X1 U295 ( .A(n24), .Z(n248) );
  BUF_X1 U296 ( .A(n18), .Z(n236) );
  BUF_X1 U297 ( .A(n25), .Z(n260) );
  BUF_X1 U298 ( .A(n44), .Z(n188) );
  BUF_X1 U299 ( .A(n41), .Z(n200) );
  BUF_X1 U300 ( .A(n16), .Z(n224) );
  BUF_X1 U301 ( .A(n45), .Z(n212) );
  BUF_X1 U302 ( .A(n26), .Z(n176) );
  AND2_X1 U303 ( .A1(n9), .A2(n11), .ZN(n5) );
  AND2_X1 U304 ( .A1(n10), .A2(n12), .ZN(n6) );
  AND2_X1 U305 ( .A1(n368), .A2(n162), .ZN(n7) );
  AND2_X1 U306 ( .A1(n368), .A2(n264), .ZN(n8) );
  AND2_X2 U307 ( .A1(n372), .A2(n371), .ZN(n9) );
  AND2_X2 U308 ( .A1(n1036), .A2(n1035), .ZN(n10) );
  BUF_X1 U309 ( .A(n1031), .Z(n163) );
  BUF_X1 U310 ( .A(n2205), .Z(n265) );
  AND2_X1 U311 ( .A1(n60), .A2(n384), .ZN(n11) );
  AND2_X1 U312 ( .A1(n61), .A2(n1058), .ZN(n12) );
  AND3_X1 U313 ( .A1(n383), .A2(n384), .A3(n374), .ZN(n13) );
  AND3_X1 U314 ( .A1(n1057), .A2(n1058), .A3(n1040), .ZN(n14) );
  CLKBUF_X1 U315 ( .A(n1031), .Z(n164) );
  CLKBUF_X1 U316 ( .A(n2205), .Z(n266) );
  AND2_X1 U317 ( .A1(n46), .A2(n48), .ZN(n15) );
  AND2_X1 U318 ( .A1(n47), .A2(n49), .ZN(n16) );
  AND2_X1 U319 ( .A1(n9), .A2(n48), .ZN(n17) );
  AND2_X1 U320 ( .A1(n10), .A2(n49), .ZN(n18) );
  AND2_X1 U321 ( .A1(n11), .A2(n46), .ZN(n19) );
  AND2_X1 U322 ( .A1(n12), .A2(n47), .ZN(n20) );
  AND2_X1 U323 ( .A1(n51), .A2(n1), .ZN(n21) );
  AND2_X1 U324 ( .A1(n51), .A2(n2), .ZN(n22) );
  AND2_X1 U325 ( .A1(n54), .A2(n1), .ZN(n23) );
  AND2_X1 U326 ( .A1(n56), .A2(n3), .ZN(n24) );
  AND2_X1 U327 ( .A1(n56), .A2(n4), .ZN(n25) );
  AND2_X1 U328 ( .A1(n58), .A2(n3), .ZN(n26) );
  AND2_X1 U329 ( .A1(n50), .A2(n1), .ZN(n27) );
  AND2_X1 U330 ( .A1(n50), .A2(n2), .ZN(n28) );
  AND2_X1 U331 ( .A1(n53), .A2(n2), .ZN(n29) );
  AND2_X1 U332 ( .A1(n13), .A2(n1), .ZN(n30) );
  AND2_X1 U333 ( .A1(n13), .A2(n2), .ZN(n31) );
  AND2_X1 U334 ( .A1(n55), .A2(n3), .ZN(n32) );
  AND2_X1 U335 ( .A1(n53), .A2(n1), .ZN(n33) );
  AND2_X1 U336 ( .A1(n55), .A2(n4), .ZN(n34) );
  AND2_X1 U337 ( .A1(n59), .A2(n4), .ZN(n35) );
  AND2_X1 U338 ( .A1(n14), .A2(n3), .ZN(n36) );
  AND2_X1 U339 ( .A1(n14), .A2(n4), .ZN(n37) );
  AND2_X1 U340 ( .A1(n59), .A2(n3), .ZN(n38) );
  INV_X1 U341 ( .A(RST), .ZN(n369) );
  AND2_X1 U342 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .ZN(n39) );
  AND2_X1 U343 ( .A1(n52), .A2(n1), .ZN(n40) );
  AND2_X1 U344 ( .A1(n57), .A2(n3), .ZN(n41) );
  AND2_X1 U345 ( .A1(n54), .A2(n2), .ZN(n42) );
  AND2_X1 U346 ( .A1(n52), .A2(n2), .ZN(n43) );
  AND2_X1 U347 ( .A1(n58), .A2(n4), .ZN(n44) );
  AND2_X1 U348 ( .A1(n57), .A2(n4), .ZN(n45) );
  AND2_X2 U349 ( .A1(ADD_RD2[2]), .A2(n372), .ZN(n46) );
  AND2_X2 U350 ( .A1(ADD_RD1[2]), .A2(n1036), .ZN(n47) );
  NAND2_X1 U351 ( .A1(DATAIN[1]), .A2(n368), .ZN(n4400) );
  NAND2_X1 U352 ( .A1(DATAIN[2]), .A2(n368), .ZN(n4402) );
  NAND2_X1 U353 ( .A1(DATAIN[3]), .A2(n368), .ZN(n4404) );
  AND2_X1 U354 ( .A1(ADD_RD2[0]), .A2(n60), .ZN(n48) );
  AND2_X1 U355 ( .A1(ADD_RD1[0]), .A2(n61), .ZN(n49) );
  AND3_X1 U356 ( .A1(ADD_RD2[4]), .A2(n384), .A3(n383), .ZN(n50) );
  AND3_X1 U357 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n383), .ZN(n51) );
  AND3_X1 U358 ( .A1(ADD_RD2[0]), .A2(n383), .A3(n374), .ZN(n52) );
  AND3_X1 U359 ( .A1(ADD_RD2[3]), .A2(n384), .A3(n374), .ZN(n53) );
  AND3_X1 U360 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n374), .ZN(n54) );
  AND3_X1 U361 ( .A1(ADD_RD1[4]), .A2(n1058), .A3(n1057), .ZN(n55) );
  AND3_X1 U362 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n1057), .ZN(n56) );
  AND3_X1 U363 ( .A1(ADD_RD1[0]), .A2(n1057), .A3(n1040), .ZN(n57) );
  AND3_X1 U364 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n1040), .ZN(n58) );
  AND3_X1 U365 ( .A1(ADD_RD1[3]), .A2(n1058), .A3(n1040), .ZN(n59) );
  AND2_X1 U366 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .ZN(n60) );
  AND2_X1 U367 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .ZN(n61) );
  AND2_X1 U368 ( .A1(ADD_WR[4]), .A2(WR), .ZN(n62) );
  INV_X1 U369 ( .A(n369), .ZN(n363) );
  INV_X1 U370 ( .A(n369), .ZN(n364) );
  INV_X1 U371 ( .A(n369), .ZN(n365) );
  INV_X1 U372 ( .A(n369), .ZN(n366) );
  INV_X1 U373 ( .A(n369), .ZN(n367) );
  INV_X1 U374 ( .A(n369), .ZN(n368) );
  OR2_X1 U375 ( .A1(RD2), .A2(n369), .ZN(n1031) );
  INV_X1 U376 ( .A(ADD_RD2[4]), .ZN(n374) );
  INV_X1 U377 ( .A(ADD_RD2[0]), .ZN(n384) );
  INV_X1 U378 ( .A(ADD_RD2[1]), .ZN(n372) );
  NAND2_X1 U379 ( .A1(n54), .A2(n46), .ZN(n996) );
  NAND2_X1 U380 ( .A1(n53), .A2(n46), .ZN(n995) );
  OAI22_X1 U381 ( .A1(n1033), .A2(n66), .B1(n1032), .B2(n63), .ZN(n370) );
  AOI221_X1 U382 ( .B1(n72), .B2(n3844), .C1(n69), .C2(n3878), .A(n370), .ZN(
        n380) );
  INV_X1 U383 ( .A(ADD_RD2[2]), .ZN(n371) );
  NAND2_X1 U384 ( .A1(n54), .A2(n9), .ZN(n999) );
  NAND2_X1 U385 ( .A1(n53), .A2(n9), .ZN(n998) );
  OAI22_X1 U386 ( .A1(n1038), .A2(n78), .B1(n1037), .B2(n75), .ZN(n373) );
  AOI221_X1 U387 ( .B1(n84), .B2(n3980), .C1(n81), .C2(n4014), .A(n373), .ZN(
        n379) );
  INV_X1 U388 ( .A(ADD_RD2[3]), .ZN(n383) );
  NAND2_X1 U389 ( .A1(n52), .A2(n46), .ZN(n1002) );
  NAND2_X1 U390 ( .A1(n13), .A2(n46), .ZN(n1001) );
  OAI22_X1 U391 ( .A1(n1042), .A2(n90), .B1(n1041), .B2(n87), .ZN(n375) );
  AOI221_X1 U392 ( .B1(n96), .B2(n4120), .C1(n93), .C2(n4155), .A(n375), .ZN(
        n378) );
  NAND2_X1 U393 ( .A1(n52), .A2(n9), .ZN(n1005) );
  NAND2_X1 U394 ( .A1(n13), .A2(n9), .ZN(n1004) );
  OAI22_X1 U395 ( .A1(n1045), .A2(n102), .B1(n1044), .B2(n99), .ZN(n376) );
  AOI221_X1 U396 ( .B1(n108), .B2(n4260), .C1(n105), .C2(n4295), .A(n376), 
        .ZN(n377) );
  NAND4_X1 U397 ( .A1(n380), .A2(n379), .A3(n378), .A4(n377), .ZN(n392) );
  NAND2_X1 U398 ( .A1(n1), .A2(n48), .ZN(n1012) );
  NAND2_X1 U399 ( .A1(n1), .A2(n11), .ZN(n1011) );
  OAI22_X1 U400 ( .A1(n1052), .A2(n114), .B1(n1051), .B2(n111), .ZN(n381) );
  AOI221_X1 U401 ( .B1(n120), .B2(n2275), .C1(n117), .C2(n2309), .A(n381), 
        .ZN(n390) );
  NAND2_X1 U402 ( .A1(n2), .A2(n48), .ZN(n1015) );
  NAND2_X1 U403 ( .A1(n2), .A2(n11), .ZN(n1014) );
  OAI22_X1 U404 ( .A1(n1055), .A2(n126), .B1(n1054), .B2(n123), .ZN(n382) );
  AOI221_X1 U405 ( .B1(n132), .B2(n2411), .C1(n129), .C2(n2449), .A(n382), 
        .ZN(n389) );
  NAND2_X1 U406 ( .A1(n51), .A2(n46), .ZN(n1018) );
  NAND2_X1 U407 ( .A1(n50), .A2(n46), .ZN(n1017) );
  OAI22_X1 U408 ( .A1(n1060), .A2(n138), .B1(n1059), .B2(n135), .ZN(n385) );
  AOI221_X1 U409 ( .B1(n144), .B2(n2483), .C1(n141), .C2(n2517), .A(n385), 
        .ZN(n388) );
  NAND2_X1 U410 ( .A1(n51), .A2(n9), .ZN(n1021) );
  NAND2_X1 U411 ( .A1(n50), .A2(n9), .ZN(n1020) );
  OAI22_X1 U412 ( .A1(n1063), .A2(n150), .B1(n1062), .B2(n147), .ZN(n386) );
  AOI221_X1 U413 ( .B1(n156), .B2(n3707), .C1(n153), .C2(n3741), .A(n386), 
        .ZN(n387) );
  NAND4_X1 U414 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(n391) );
  OAI21_X1 U415 ( .B1(n392), .B2(n391), .A(n159), .ZN(n393) );
  OAI21_X1 U416 ( .B1(n162), .B2(n394), .A(n393), .ZN(n2527) );
  OAI22_X1 U417 ( .A1(n1074), .A2(n66), .B1(n1073), .B2(n63), .ZN(n395) );
  AOI221_X1 U418 ( .B1(n72), .B2(n3845), .C1(n69), .C2(n3879), .A(n395), .ZN(
        n402) );
  OAI22_X1 U419 ( .A1(n1077), .A2(n78), .B1(n1076), .B2(n75), .ZN(n396) );
  AOI221_X1 U420 ( .B1(n84), .B2(n3981), .C1(n81), .C2(n4015), .A(n396), .ZN(
        n401) );
  OAI22_X1 U421 ( .A1(n1080), .A2(n90), .B1(n1079), .B2(n87), .ZN(n397) );
  AOI221_X1 U422 ( .B1(n96), .B2(n4121), .C1(n93), .C2(n4156), .A(n397), .ZN(
        n400) );
  OAI22_X1 U423 ( .A1(n1083), .A2(n102), .B1(n1082), .B2(n99), .ZN(n398) );
  AOI221_X1 U424 ( .B1(n108), .B2(n4261), .C1(n105), .C2(n4297), .A(n398), 
        .ZN(n399) );
  NAND4_X1 U425 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(n412) );
  OAI22_X1 U426 ( .A1(n1090), .A2(n114), .B1(n1089), .B2(n111), .ZN(n403) );
  AOI221_X1 U427 ( .B1(n120), .B2(n2276), .C1(n117), .C2(n2310), .A(n403), 
        .ZN(n410) );
  OAI22_X1 U428 ( .A1(n1093), .A2(n126), .B1(n1092), .B2(n123), .ZN(n404) );
  AOI221_X1 U429 ( .B1(n132), .B2(n2412), .C1(n129), .C2(n2450), .A(n404), 
        .ZN(n409) );
  OAI22_X1 U430 ( .A1(n1096), .A2(n138), .B1(n1095), .B2(n135), .ZN(n405) );
  AOI221_X1 U431 ( .B1(n144), .B2(n2484), .C1(n141), .C2(n2518), .A(n405), 
        .ZN(n408) );
  OAI22_X1 U432 ( .A1(n1099), .A2(n150), .B1(n1098), .B2(n147), .ZN(n406) );
  AOI221_X1 U433 ( .B1(n156), .B2(n3708), .C1(n153), .C2(n3742), .A(n406), 
        .ZN(n407) );
  NAND4_X1 U434 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(n411) );
  OAI21_X1 U435 ( .B1(n412), .B2(n411), .A(n159), .ZN(n413) );
  OAI21_X1 U436 ( .B1(n162), .B2(n414), .A(n413), .ZN(n2528) );
  OAI22_X1 U437 ( .A1(n1110), .A2(n66), .B1(n1109), .B2(n63), .ZN(n415) );
  AOI221_X1 U438 ( .B1(n72), .B2(n3846), .C1(n69), .C2(n3880), .A(n415), .ZN(
        n422) );
  OAI22_X1 U439 ( .A1(n1113), .A2(n78), .B1(n1112), .B2(n75), .ZN(n416) );
  AOI221_X1 U440 ( .B1(n84), .B2(n3982), .C1(n81), .C2(n4016), .A(n416), .ZN(
        n421) );
  OAI22_X1 U441 ( .A1(n1116), .A2(n90), .B1(n1115), .B2(n87), .ZN(n417) );
  AOI221_X1 U442 ( .B1(n96), .B2(n4122), .C1(n93), .C2(n4157), .A(n417), .ZN(
        n420) );
  OAI22_X1 U443 ( .A1(n1119), .A2(n102), .B1(n1118), .B2(n99), .ZN(n418) );
  AOI221_X1 U444 ( .B1(n108), .B2(n4262), .C1(n105), .C2(n4299), .A(n418), 
        .ZN(n419) );
  NAND4_X1 U445 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(n432) );
  OAI22_X1 U446 ( .A1(n1126), .A2(n114), .B1(n1125), .B2(n111), .ZN(n423) );
  AOI221_X1 U447 ( .B1(n120), .B2(n2277), .C1(n117), .C2(n2311), .A(n423), 
        .ZN(n430) );
  OAI22_X1 U448 ( .A1(n1129), .A2(n126), .B1(n1128), .B2(n123), .ZN(n424) );
  AOI221_X1 U449 ( .B1(n132), .B2(n2413), .C1(n129), .C2(n2451), .A(n424), 
        .ZN(n429) );
  OAI22_X1 U450 ( .A1(n1132), .A2(n138), .B1(n1131), .B2(n135), .ZN(n425) );
  AOI221_X1 U451 ( .B1(n144), .B2(n2485), .C1(n141), .C2(n2519), .A(n425), 
        .ZN(n428) );
  OAI22_X1 U452 ( .A1(n1135), .A2(n150), .B1(n1134), .B2(n147), .ZN(n426) );
  AOI221_X1 U453 ( .B1(n156), .B2(n3709), .C1(n153), .C2(n3743), .A(n426), 
        .ZN(n427) );
  NAND4_X1 U454 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(n431) );
  OAI21_X1 U455 ( .B1(n432), .B2(n431), .A(n159), .ZN(n433) );
  OAI21_X1 U456 ( .B1(n162), .B2(n434), .A(n433), .ZN(n2529) );
  OAI22_X1 U457 ( .A1(n1146), .A2(n66), .B1(n1145), .B2(n63), .ZN(n435) );
  AOI221_X1 U458 ( .B1(n72), .B2(n3847), .C1(n69), .C2(n3881), .A(n435), .ZN(
        n442) );
  OAI22_X1 U459 ( .A1(n1149), .A2(n78), .B1(n1148), .B2(n75), .ZN(n436) );
  AOI221_X1 U460 ( .B1(n84), .B2(n3983), .C1(n81), .C2(n4017), .A(n436), .ZN(
        n441) );
  OAI22_X1 U461 ( .A1(n1152), .A2(n90), .B1(n1151), .B2(n87), .ZN(n437) );
  AOI221_X1 U462 ( .B1(n96), .B2(n4123), .C1(n93), .C2(n4158), .A(n437), .ZN(
        n440) );
  OAI22_X1 U463 ( .A1(n1155), .A2(n102), .B1(n1154), .B2(n99), .ZN(n438) );
  AOI221_X1 U464 ( .B1(n108), .B2(n4263), .C1(n105), .C2(n4301), .A(n438), 
        .ZN(n439) );
  NAND4_X1 U465 ( .A1(n442), .A2(n441), .A3(n440), .A4(n439), .ZN(n452) );
  OAI22_X1 U466 ( .A1(n1162), .A2(n114), .B1(n1161), .B2(n111), .ZN(n443) );
  AOI221_X1 U467 ( .B1(n120), .B2(n2278), .C1(n117), .C2(n2312), .A(n443), 
        .ZN(n450) );
  OAI22_X1 U468 ( .A1(n1165), .A2(n126), .B1(n1164), .B2(n123), .ZN(n444) );
  AOI221_X1 U469 ( .B1(n132), .B2(n2414), .C1(n129), .C2(n2452), .A(n444), 
        .ZN(n449) );
  OAI22_X1 U470 ( .A1(n1168), .A2(n138), .B1(n1167), .B2(n135), .ZN(n445) );
  AOI221_X1 U471 ( .B1(n144), .B2(n2486), .C1(n141), .C2(n2520), .A(n445), 
        .ZN(n448) );
  OAI22_X1 U472 ( .A1(n1171), .A2(n150), .B1(n1170), .B2(n147), .ZN(n446) );
  AOI221_X1 U473 ( .B1(n156), .B2(n3710), .C1(n153), .C2(n3744), .A(n446), 
        .ZN(n447) );
  NAND4_X1 U474 ( .A1(n450), .A2(n449), .A3(n448), .A4(n447), .ZN(n451) );
  OAI21_X1 U475 ( .B1(n452), .B2(n451), .A(n159), .ZN(n453) );
  OAI21_X1 U476 ( .B1(n162), .B2(n454), .A(n453), .ZN(n2530) );
  OAI22_X1 U477 ( .A1(n1182), .A2(n66), .B1(n1181), .B2(n63), .ZN(n455) );
  AOI221_X1 U478 ( .B1(n72), .B2(n3848), .C1(n69), .C2(n3882), .A(n455), .ZN(
        n462) );
  OAI22_X1 U479 ( .A1(n1185), .A2(n78), .B1(n1184), .B2(n75), .ZN(n456) );
  AOI221_X1 U480 ( .B1(n84), .B2(n3984), .C1(n81), .C2(n4018), .A(n456), .ZN(
        n461) );
  OAI22_X1 U481 ( .A1(n1188), .A2(n90), .B1(n1187), .B2(n87), .ZN(n457) );
  AOI221_X1 U482 ( .B1(n96), .B2(n4124), .C1(n93), .C2(n4159), .A(n457), .ZN(
        n460) );
  OAI22_X1 U483 ( .A1(n1191), .A2(n102), .B1(n1190), .B2(n99), .ZN(n458) );
  AOI221_X1 U484 ( .B1(n108), .B2(n4264), .C1(n105), .C2(n4303), .A(n458), 
        .ZN(n459) );
  NAND4_X1 U485 ( .A1(n462), .A2(n461), .A3(n460), .A4(n459), .ZN(n472) );
  OAI22_X1 U486 ( .A1(n1198), .A2(n114), .B1(n1197), .B2(n111), .ZN(n463) );
  AOI221_X1 U487 ( .B1(n120), .B2(n2279), .C1(n117), .C2(n2313), .A(n463), 
        .ZN(n470) );
  OAI22_X1 U488 ( .A1(n1201), .A2(n126), .B1(n1200), .B2(n123), .ZN(n464) );
  AOI221_X1 U489 ( .B1(n132), .B2(n2415), .C1(n129), .C2(n2453), .A(n464), 
        .ZN(n469) );
  OAI22_X1 U490 ( .A1(n1204), .A2(n138), .B1(n1203), .B2(n135), .ZN(n465) );
  AOI221_X1 U491 ( .B1(n144), .B2(n2487), .C1(n141), .C2(n2521), .A(n465), 
        .ZN(n468) );
  OAI22_X1 U492 ( .A1(n1207), .A2(n150), .B1(n1206), .B2(n147), .ZN(n466) );
  AOI221_X1 U493 ( .B1(n156), .B2(n3711), .C1(n153), .C2(n3745), .A(n466), 
        .ZN(n467) );
  NAND4_X1 U494 ( .A1(n470), .A2(n469), .A3(n468), .A4(n467), .ZN(n471) );
  OAI21_X1 U495 ( .B1(n472), .B2(n471), .A(n159), .ZN(n473) );
  OAI21_X1 U496 ( .B1(n162), .B2(n474), .A(n473), .ZN(n2531) );
  OAI22_X1 U497 ( .A1(n1218), .A2(n66), .B1(n1217), .B2(n63), .ZN(n475) );
  AOI221_X1 U498 ( .B1(n72), .B2(n3849), .C1(n69), .C2(n3883), .A(n475), .ZN(
        n482) );
  OAI22_X1 U499 ( .A1(n1221), .A2(n78), .B1(n1220), .B2(n75), .ZN(n476) );
  AOI221_X1 U500 ( .B1(n84), .B2(n3985), .C1(n81), .C2(n4019), .A(n476), .ZN(
        n481) );
  OAI22_X1 U501 ( .A1(n1224), .A2(n90), .B1(n1223), .B2(n87), .ZN(n477) );
  AOI221_X1 U502 ( .B1(n96), .B2(n4125), .C1(n93), .C2(n4160), .A(n477), .ZN(
        n480) );
  OAI22_X1 U503 ( .A1(n1227), .A2(n102), .B1(n1226), .B2(n99), .ZN(n478) );
  AOI221_X1 U504 ( .B1(n108), .B2(n4265), .C1(n105), .C2(n4305), .A(n478), 
        .ZN(n479) );
  NAND4_X1 U505 ( .A1(n482), .A2(n481), .A3(n480), .A4(n479), .ZN(n492) );
  OAI22_X1 U506 ( .A1(n1234), .A2(n114), .B1(n1233), .B2(n111), .ZN(n483) );
  AOI221_X1 U507 ( .B1(n120), .B2(n2280), .C1(n117), .C2(n2314), .A(n483), 
        .ZN(n490) );
  OAI22_X1 U508 ( .A1(n1237), .A2(n126), .B1(n1236), .B2(n123), .ZN(n484) );
  AOI221_X1 U509 ( .B1(n132), .B2(n2416), .C1(n129), .C2(n2454), .A(n484), 
        .ZN(n489) );
  OAI22_X1 U510 ( .A1(n1240), .A2(n138), .B1(n1239), .B2(n135), .ZN(n485) );
  AOI221_X1 U511 ( .B1(n144), .B2(n2488), .C1(n141), .C2(n2522), .A(n485), 
        .ZN(n488) );
  OAI22_X1 U512 ( .A1(n1243), .A2(n150), .B1(n1242), .B2(n147), .ZN(n486) );
  AOI221_X1 U513 ( .B1(n156), .B2(n3712), .C1(n153), .C2(n3746), .A(n486), 
        .ZN(n487) );
  NAND4_X1 U514 ( .A1(n490), .A2(n489), .A3(n488), .A4(n487), .ZN(n491) );
  OAI21_X1 U515 ( .B1(n492), .B2(n491), .A(n159), .ZN(n493) );
  OAI21_X1 U516 ( .B1(n162), .B2(n494), .A(n493), .ZN(n2532) );
  OAI22_X1 U517 ( .A1(n1254), .A2(n66), .B1(n1253), .B2(n63), .ZN(n495) );
  AOI221_X1 U518 ( .B1(n72), .B2(n3850), .C1(n69), .C2(n3884), .A(n495), .ZN(
        n502) );
  OAI22_X1 U519 ( .A1(n1257), .A2(n78), .B1(n1256), .B2(n75), .ZN(n496) );
  AOI221_X1 U520 ( .B1(n84), .B2(n3986), .C1(n81), .C2(n4020), .A(n496), .ZN(
        n501) );
  OAI22_X1 U521 ( .A1(n1260), .A2(n90), .B1(n1259), .B2(n87), .ZN(n497) );
  AOI221_X1 U522 ( .B1(n96), .B2(n4126), .C1(n93), .C2(n4161), .A(n497), .ZN(
        n500) );
  OAI22_X1 U523 ( .A1(n1263), .A2(n102), .B1(n1262), .B2(n99), .ZN(n498) );
  AOI221_X1 U524 ( .B1(n108), .B2(n4266), .C1(n105), .C2(n4307), .A(n498), 
        .ZN(n499) );
  NAND4_X1 U525 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .ZN(n512) );
  OAI22_X1 U526 ( .A1(n1270), .A2(n114), .B1(n1269), .B2(n111), .ZN(n503) );
  AOI221_X1 U527 ( .B1(n120), .B2(n2281), .C1(n117), .C2(n2315), .A(n503), 
        .ZN(n510) );
  OAI22_X1 U528 ( .A1(n1273), .A2(n126), .B1(n1272), .B2(n123), .ZN(n504) );
  AOI221_X1 U529 ( .B1(n132), .B2(n2417), .C1(n129), .C2(n2455), .A(n504), 
        .ZN(n509) );
  OAI22_X1 U530 ( .A1(n1276), .A2(n138), .B1(n1275), .B2(n135), .ZN(n505) );
  AOI221_X1 U531 ( .B1(n144), .B2(n2489), .C1(n141), .C2(n2523), .A(n505), 
        .ZN(n508) );
  OAI22_X1 U532 ( .A1(n1279), .A2(n150), .B1(n1278), .B2(n147), .ZN(n506) );
  AOI221_X1 U533 ( .B1(n156), .B2(n3713), .C1(n153), .C2(n3747), .A(n506), 
        .ZN(n507) );
  NAND4_X1 U534 ( .A1(n510), .A2(n509), .A3(n508), .A4(n507), .ZN(n511) );
  OAI21_X1 U535 ( .B1(n512), .B2(n511), .A(n159), .ZN(n513) );
  OAI21_X1 U536 ( .B1(n162), .B2(n514), .A(n513), .ZN(n2533) );
  OAI22_X1 U537 ( .A1(n1290), .A2(n66), .B1(n1289), .B2(n63), .ZN(n515) );
  AOI221_X1 U538 ( .B1(n72), .B2(n3851), .C1(n69), .C2(n3885), .A(n515), .ZN(
        n522) );
  OAI22_X1 U539 ( .A1(n1293), .A2(n78), .B1(n1292), .B2(n75), .ZN(n516) );
  AOI221_X1 U540 ( .B1(n84), .B2(n3987), .C1(n81), .C2(n4021), .A(n516), .ZN(
        n521) );
  OAI22_X1 U541 ( .A1(n1296), .A2(n90), .B1(n1295), .B2(n87), .ZN(n517) );
  AOI221_X1 U542 ( .B1(n96), .B2(n4127), .C1(n93), .C2(n4162), .A(n517), .ZN(
        n520) );
  OAI22_X1 U543 ( .A1(n1299), .A2(n102), .B1(n1298), .B2(n99), .ZN(n518) );
  AOI221_X1 U544 ( .B1(n108), .B2(n4267), .C1(n105), .C2(n4309), .A(n518), 
        .ZN(n519) );
  NAND4_X1 U545 ( .A1(n522), .A2(n521), .A3(n520), .A4(n519), .ZN(n532) );
  OAI22_X1 U546 ( .A1(n1306), .A2(n114), .B1(n1305), .B2(n111), .ZN(n523) );
  AOI221_X1 U547 ( .B1(n120), .B2(n2282), .C1(n117), .C2(n2316), .A(n523), 
        .ZN(n530) );
  OAI22_X1 U548 ( .A1(n1309), .A2(n126), .B1(n1308), .B2(n123), .ZN(n524) );
  AOI221_X1 U549 ( .B1(n132), .B2(n2418), .C1(n129), .C2(n2456), .A(n524), 
        .ZN(n529) );
  OAI22_X1 U550 ( .A1(n1312), .A2(n138), .B1(n1311), .B2(n135), .ZN(n525) );
  AOI221_X1 U551 ( .B1(n144), .B2(n2490), .C1(n141), .C2(n2524), .A(n525), 
        .ZN(n528) );
  OAI22_X1 U552 ( .A1(n1315), .A2(n150), .B1(n1314), .B2(n147), .ZN(n526) );
  AOI221_X1 U553 ( .B1(n156), .B2(n3714), .C1(n153), .C2(n3748), .A(n526), 
        .ZN(n527) );
  NAND4_X1 U554 ( .A1(n530), .A2(n529), .A3(n528), .A4(n527), .ZN(n531) );
  OAI21_X1 U555 ( .B1(n532), .B2(n531), .A(n159), .ZN(n533) );
  OAI21_X1 U556 ( .B1(n162), .B2(n534), .A(n533), .ZN(n2534) );
  OAI22_X1 U557 ( .A1(n1326), .A2(n66), .B1(n1325), .B2(n63), .ZN(n535) );
  AOI221_X1 U558 ( .B1(n72), .B2(n3852), .C1(n69), .C2(n3886), .A(n535), .ZN(
        n542) );
  OAI22_X1 U559 ( .A1(n1329), .A2(n78), .B1(n1328), .B2(n75), .ZN(n536) );
  AOI221_X1 U560 ( .B1(n84), .B2(n3988), .C1(n81), .C2(n4022), .A(n536), .ZN(
        n541) );
  OAI22_X1 U561 ( .A1(n1332), .A2(n90), .B1(n1331), .B2(n87), .ZN(n537) );
  AOI221_X1 U562 ( .B1(n96), .B2(n4128), .C1(n93), .C2(n4163), .A(n537), .ZN(
        n540) );
  OAI22_X1 U563 ( .A1(n1335), .A2(n102), .B1(n1334), .B2(n99), .ZN(n538) );
  AOI221_X1 U564 ( .B1(n108), .B2(n4268), .C1(n105), .C2(n4311), .A(n538), 
        .ZN(n539) );
  NAND4_X1 U565 ( .A1(n542), .A2(n541), .A3(n540), .A4(n539), .ZN(n552) );
  OAI22_X1 U566 ( .A1(n1342), .A2(n114), .B1(n1341), .B2(n111), .ZN(n543) );
  AOI221_X1 U567 ( .B1(n120), .B2(n2283), .C1(n117), .C2(n2317), .A(n543), 
        .ZN(n550) );
  OAI22_X1 U568 ( .A1(n1345), .A2(n126), .B1(n1344), .B2(n123), .ZN(n544) );
  AOI221_X1 U569 ( .B1(n132), .B2(n2419), .C1(n129), .C2(n2457), .A(n544), 
        .ZN(n549) );
  OAI22_X1 U570 ( .A1(n1348), .A2(n138), .B1(n1347), .B2(n135), .ZN(n545) );
  AOI221_X1 U571 ( .B1(n144), .B2(n2491), .C1(n141), .C2(n2525), .A(n545), 
        .ZN(n548) );
  OAI22_X1 U572 ( .A1(n1351), .A2(n150), .B1(n1350), .B2(n147), .ZN(n546) );
  AOI221_X1 U573 ( .B1(n156), .B2(n3715), .C1(n153), .C2(n3749), .A(n546), 
        .ZN(n547) );
  NAND4_X1 U574 ( .A1(n550), .A2(n549), .A3(n548), .A4(n547), .ZN(n551) );
  OAI21_X1 U575 ( .B1(n552), .B2(n551), .A(n159), .ZN(n553) );
  OAI21_X1 U576 ( .B1(n162), .B2(n554), .A(n553), .ZN(n2535) );
  OAI22_X1 U577 ( .A1(n1362), .A2(n66), .B1(n1361), .B2(n63), .ZN(n555) );
  AOI221_X1 U578 ( .B1(n72), .B2(n3853), .C1(n69), .C2(n3887), .A(n555), .ZN(
        n562) );
  OAI22_X1 U579 ( .A1(n1365), .A2(n78), .B1(n1364), .B2(n75), .ZN(n556) );
  AOI221_X1 U580 ( .B1(n84), .B2(n3989), .C1(n81), .C2(n4023), .A(n556), .ZN(
        n561) );
  OAI22_X1 U581 ( .A1(n1368), .A2(n90), .B1(n1367), .B2(n87), .ZN(n557) );
  AOI221_X1 U582 ( .B1(n96), .B2(n4129), .C1(n93), .C2(n4164), .A(n557), .ZN(
        n560) );
  OAI22_X1 U583 ( .A1(n1371), .A2(n102), .B1(n1370), .B2(n99), .ZN(n558) );
  AOI221_X1 U584 ( .B1(n108), .B2(n4269), .C1(n105), .C2(n4313), .A(n558), 
        .ZN(n559) );
  NAND4_X1 U585 ( .A1(n562), .A2(n561), .A3(n560), .A4(n559), .ZN(n572) );
  OAI22_X1 U586 ( .A1(n1378), .A2(n114), .B1(n1377), .B2(n111), .ZN(n563) );
  AOI221_X1 U587 ( .B1(n120), .B2(n2284), .C1(n117), .C2(n2318), .A(n563), 
        .ZN(n570) );
  OAI22_X1 U588 ( .A1(n1381), .A2(n126), .B1(n1380), .B2(n123), .ZN(n564) );
  AOI221_X1 U589 ( .B1(n132), .B2(n2420), .C1(n129), .C2(n2458), .A(n564), 
        .ZN(n569) );
  OAI22_X1 U590 ( .A1(n1384), .A2(n138), .B1(n1383), .B2(n135), .ZN(n565) );
  AOI221_X1 U591 ( .B1(n144), .B2(n2492), .C1(n141), .C2(n2526), .A(n565), 
        .ZN(n568) );
  OAI22_X1 U592 ( .A1(n1387), .A2(n150), .B1(n1386), .B2(n147), .ZN(n566) );
  AOI221_X1 U593 ( .B1(n156), .B2(n3716), .C1(n153), .C2(n3750), .A(n566), 
        .ZN(n567) );
  NAND4_X1 U594 ( .A1(n570), .A2(n569), .A3(n568), .A4(n567), .ZN(n571) );
  OAI21_X1 U595 ( .B1(n572), .B2(n571), .A(n159), .ZN(n573) );
  OAI21_X1 U596 ( .B1(n162), .B2(n574), .A(n573), .ZN(n2536) );
  OAI22_X1 U597 ( .A1(n1398), .A2(n66), .B1(n1397), .B2(n63), .ZN(n575) );
  AOI221_X1 U598 ( .B1(n72), .B2(n3854), .C1(n69), .C2(n3888), .A(n575), .ZN(
        n582) );
  OAI22_X1 U599 ( .A1(n1401), .A2(n78), .B1(n1400), .B2(n75), .ZN(n576) );
  AOI221_X1 U600 ( .B1(n84), .B2(n3990), .C1(n81), .C2(n4024), .A(n576), .ZN(
        n581) );
  OAI22_X1 U601 ( .A1(n1404), .A2(n90), .B1(n1403), .B2(n87), .ZN(n577) );
  AOI221_X1 U602 ( .B1(n96), .B2(n4130), .C1(n93), .C2(n4165), .A(n577), .ZN(
        n580) );
  OAI22_X1 U603 ( .A1(n1407), .A2(n102), .B1(n1406), .B2(n99), .ZN(n578) );
  AOI221_X1 U604 ( .B1(n108), .B2(n4270), .C1(n105), .C2(n4315), .A(n578), 
        .ZN(n579) );
  NAND4_X1 U605 ( .A1(n582), .A2(n581), .A3(n580), .A4(n579), .ZN(n592) );
  OAI22_X1 U606 ( .A1(n1414), .A2(n114), .B1(n1413), .B2(n111), .ZN(n583) );
  AOI221_X1 U607 ( .B1(n120), .B2(n2285), .C1(n117), .C2(n2319), .A(n583), 
        .ZN(n590) );
  OAI22_X1 U608 ( .A1(n1417), .A2(n126), .B1(n1416), .B2(n123), .ZN(n584) );
  AOI221_X1 U609 ( .B1(n132), .B2(n2421), .C1(n129), .C2(n2459), .A(n584), 
        .ZN(n589) );
  OAI22_X1 U610 ( .A1(n1420), .A2(n138), .B1(n1419), .B2(n135), .ZN(n585) );
  AOI221_X1 U611 ( .B1(n144), .B2(n2493), .C1(n141), .C2(n3615), .A(n585), 
        .ZN(n588) );
  OAI22_X1 U612 ( .A1(n1423), .A2(n150), .B1(n1422), .B2(n147), .ZN(n586) );
  AOI221_X1 U613 ( .B1(n156), .B2(n3717), .C1(n153), .C2(n3751), .A(n586), 
        .ZN(n587) );
  NAND4_X1 U614 ( .A1(n590), .A2(n589), .A3(n588), .A4(n587), .ZN(n591) );
  OAI21_X1 U615 ( .B1(n592), .B2(n591), .A(n159), .ZN(n593) );
  OAI21_X1 U616 ( .B1(n162), .B2(n594), .A(n593), .ZN(n2537) );
  OAI22_X1 U617 ( .A1(n1434), .A2(n66), .B1(n1433), .B2(n63), .ZN(n595) );
  AOI221_X1 U618 ( .B1(n72), .B2(n3855), .C1(n69), .C2(n3889), .A(n595), .ZN(
        n602) );
  OAI22_X1 U619 ( .A1(n1437), .A2(n78), .B1(n1436), .B2(n75), .ZN(n596) );
  AOI221_X1 U620 ( .B1(n84), .B2(n3991), .C1(n81), .C2(n4025), .A(n596), .ZN(
        n601) );
  OAI22_X1 U621 ( .A1(n1440), .A2(n90), .B1(n1439), .B2(n87), .ZN(n597) );
  AOI221_X1 U622 ( .B1(n96), .B2(n4131), .C1(n93), .C2(n4166), .A(n597), .ZN(
        n600) );
  OAI22_X1 U623 ( .A1(n1443), .A2(n102), .B1(n1442), .B2(n99), .ZN(n598) );
  AOI221_X1 U624 ( .B1(n108), .B2(n4271), .C1(n105), .C2(n4317), .A(n598), 
        .ZN(n599) );
  NAND4_X1 U625 ( .A1(n602), .A2(n601), .A3(n600), .A4(n599), .ZN(n612) );
  OAI22_X1 U626 ( .A1(n1450), .A2(n114), .B1(n1449), .B2(n111), .ZN(n603) );
  AOI221_X1 U627 ( .B1(n120), .B2(n2286), .C1(n117), .C2(n2320), .A(n603), 
        .ZN(n610) );
  OAI22_X1 U628 ( .A1(n1453), .A2(n126), .B1(n1452), .B2(n123), .ZN(n604) );
  AOI221_X1 U629 ( .B1(n132), .B2(n2422), .C1(n129), .C2(n2460), .A(n604), 
        .ZN(n609) );
  OAI22_X1 U630 ( .A1(n1456), .A2(n138), .B1(n1455), .B2(n135), .ZN(n605) );
  AOI221_X1 U631 ( .B1(n144), .B2(n2494), .C1(n141), .C2(n3616), .A(n605), 
        .ZN(n608) );
  OAI22_X1 U632 ( .A1(n1459), .A2(n150), .B1(n1458), .B2(n147), .ZN(n606) );
  AOI221_X1 U633 ( .B1(n156), .B2(n3718), .C1(n153), .C2(n3752), .A(n606), 
        .ZN(n607) );
  NAND4_X1 U634 ( .A1(n610), .A2(n609), .A3(n608), .A4(n607), .ZN(n611) );
  OAI21_X1 U635 ( .B1(n612), .B2(n611), .A(n159), .ZN(n613) );
  OAI21_X1 U636 ( .B1(n163), .B2(n614), .A(n613), .ZN(n2538) );
  OAI22_X1 U637 ( .A1(n1470), .A2(n67), .B1(n1469), .B2(n64), .ZN(n615) );
  AOI221_X1 U638 ( .B1(n73), .B2(n3856), .C1(n70), .C2(n3890), .A(n615), .ZN(
        n622) );
  OAI22_X1 U639 ( .A1(n1473), .A2(n79), .B1(n1472), .B2(n76), .ZN(n616) );
  AOI221_X1 U640 ( .B1(n85), .B2(n3992), .C1(n82), .C2(n4026), .A(n616), .ZN(
        n621) );
  OAI22_X1 U641 ( .A1(n1476), .A2(n91), .B1(n1475), .B2(n88), .ZN(n617) );
  AOI221_X1 U642 ( .B1(n97), .B2(n4132), .C1(n94), .C2(n4167), .A(n617), .ZN(
        n620) );
  OAI22_X1 U643 ( .A1(n1479), .A2(n103), .B1(n1478), .B2(n100), .ZN(n618) );
  AOI221_X1 U644 ( .B1(n109), .B2(n4272), .C1(n106), .C2(n4319), .A(n618), 
        .ZN(n619) );
  NAND4_X1 U645 ( .A1(n622), .A2(n621), .A3(n620), .A4(n619), .ZN(n632) );
  OAI22_X1 U646 ( .A1(n1486), .A2(n115), .B1(n1485), .B2(n112), .ZN(n623) );
  AOI221_X1 U647 ( .B1(n121), .B2(n2287), .C1(n118), .C2(n2321), .A(n623), 
        .ZN(n630) );
  OAI22_X1 U648 ( .A1(n1489), .A2(n127), .B1(n1488), .B2(n124), .ZN(n624) );
  AOI221_X1 U649 ( .B1(n133), .B2(n2423), .C1(n130), .C2(n2461), .A(n624), 
        .ZN(n629) );
  OAI22_X1 U650 ( .A1(n1492), .A2(n139), .B1(n1491), .B2(n136), .ZN(n625) );
  AOI221_X1 U651 ( .B1(n145), .B2(n2495), .C1(n142), .C2(n3617), .A(n625), 
        .ZN(n628) );
  OAI22_X1 U652 ( .A1(n1495), .A2(n151), .B1(n1494), .B2(n148), .ZN(n626) );
  AOI221_X1 U653 ( .B1(n157), .B2(n3719), .C1(n154), .C2(n3753), .A(n626), 
        .ZN(n627) );
  NAND4_X1 U654 ( .A1(n630), .A2(n629), .A3(n628), .A4(n627), .ZN(n631) );
  OAI21_X1 U655 ( .B1(n632), .B2(n631), .A(n160), .ZN(n633) );
  OAI21_X1 U656 ( .B1(n163), .B2(n634), .A(n633), .ZN(n2539) );
  OAI22_X1 U657 ( .A1(n1506), .A2(n67), .B1(n1505), .B2(n64), .ZN(n635) );
  AOI221_X1 U658 ( .B1(n73), .B2(n3857), .C1(n70), .C2(n3891), .A(n635), .ZN(
        n642) );
  OAI22_X1 U659 ( .A1(n1509), .A2(n79), .B1(n1508), .B2(n76), .ZN(n636) );
  AOI221_X1 U660 ( .B1(n85), .B2(n3993), .C1(n82), .C2(n4027), .A(n636), .ZN(
        n641) );
  OAI22_X1 U661 ( .A1(n1512), .A2(n91), .B1(n1511), .B2(n88), .ZN(n637) );
  AOI221_X1 U662 ( .B1(n97), .B2(n4133), .C1(n94), .C2(n4168), .A(n637), .ZN(
        n640) );
  OAI22_X1 U663 ( .A1(n1515), .A2(n103), .B1(n1514), .B2(n100), .ZN(n638) );
  AOI221_X1 U664 ( .B1(n109), .B2(n4273), .C1(n106), .C2(n4321), .A(n638), 
        .ZN(n639) );
  NAND4_X1 U665 ( .A1(n642), .A2(n641), .A3(n640), .A4(n639), .ZN(n652) );
  OAI22_X1 U666 ( .A1(n1522), .A2(n115), .B1(n1521), .B2(n112), .ZN(n643) );
  AOI221_X1 U667 ( .B1(n121), .B2(n2288), .C1(n118), .C2(n2322), .A(n643), 
        .ZN(n650) );
  OAI22_X1 U668 ( .A1(n1525), .A2(n127), .B1(n1524), .B2(n124), .ZN(n644) );
  AOI221_X1 U669 ( .B1(n133), .B2(n2424), .C1(n130), .C2(n2462), .A(n644), 
        .ZN(n649) );
  OAI22_X1 U670 ( .A1(n1528), .A2(n139), .B1(n1527), .B2(n136), .ZN(n645) );
  AOI221_X1 U671 ( .B1(n145), .B2(n2496), .C1(n142), .C2(n3618), .A(n645), 
        .ZN(n648) );
  OAI22_X1 U672 ( .A1(n1531), .A2(n151), .B1(n1530), .B2(n148), .ZN(n646) );
  AOI221_X1 U673 ( .B1(n157), .B2(n3720), .C1(n154), .C2(n3754), .A(n646), 
        .ZN(n647) );
  NAND4_X1 U674 ( .A1(n650), .A2(n649), .A3(n648), .A4(n647), .ZN(n651) );
  OAI21_X1 U675 ( .B1(n652), .B2(n651), .A(n160), .ZN(n653) );
  OAI21_X1 U676 ( .B1(n163), .B2(n654), .A(n653), .ZN(n2540) );
  OAI22_X1 U677 ( .A1(n1542), .A2(n67), .B1(n1541), .B2(n64), .ZN(n655) );
  AOI221_X1 U678 ( .B1(n73), .B2(n3858), .C1(n70), .C2(n3892), .A(n655), .ZN(
        n662) );
  OAI22_X1 U679 ( .A1(n1545), .A2(n79), .B1(n1544), .B2(n76), .ZN(n656) );
  AOI221_X1 U680 ( .B1(n85), .B2(n3994), .C1(n82), .C2(n4028), .A(n656), .ZN(
        n661) );
  OAI22_X1 U681 ( .A1(n1548), .A2(n91), .B1(n1547), .B2(n88), .ZN(n657) );
  AOI221_X1 U682 ( .B1(n97), .B2(n4134), .C1(n94), .C2(n4169), .A(n657), .ZN(
        n660) );
  OAI22_X1 U683 ( .A1(n1551), .A2(n103), .B1(n1550), .B2(n100), .ZN(n658) );
  AOI221_X1 U684 ( .B1(n109), .B2(n4274), .C1(n106), .C2(n4323), .A(n658), 
        .ZN(n659) );
  NAND4_X1 U685 ( .A1(n662), .A2(n661), .A3(n660), .A4(n659), .ZN(n672) );
  OAI22_X1 U686 ( .A1(n1558), .A2(n115), .B1(n1557), .B2(n112), .ZN(n663) );
  AOI221_X1 U687 ( .B1(n121), .B2(n2289), .C1(n118), .C2(n2323), .A(n663), 
        .ZN(n670) );
  OAI22_X1 U688 ( .A1(n1561), .A2(n127), .B1(n1560), .B2(n124), .ZN(n664) );
  AOI221_X1 U689 ( .B1(n133), .B2(n2425), .C1(n130), .C2(n2463), .A(n664), 
        .ZN(n669) );
  OAI22_X1 U690 ( .A1(n1564), .A2(n139), .B1(n1563), .B2(n136), .ZN(n665) );
  AOI221_X1 U691 ( .B1(n145), .B2(n2497), .C1(n142), .C2(n3619), .A(n665), 
        .ZN(n668) );
  OAI22_X1 U692 ( .A1(n1567), .A2(n151), .B1(n1566), .B2(n148), .ZN(n666) );
  AOI221_X1 U693 ( .B1(n157), .B2(n3721), .C1(n154), .C2(n3755), .A(n666), 
        .ZN(n667) );
  NAND4_X1 U694 ( .A1(n670), .A2(n669), .A3(n668), .A4(n667), .ZN(n671) );
  OAI21_X1 U695 ( .B1(n672), .B2(n671), .A(n160), .ZN(n673) );
  OAI21_X1 U696 ( .B1(n163), .B2(n674), .A(n673), .ZN(n2541) );
  OAI22_X1 U697 ( .A1(n1578), .A2(n67), .B1(n1577), .B2(n64), .ZN(n675) );
  AOI221_X1 U698 ( .B1(n73), .B2(n3859), .C1(n70), .C2(n3893), .A(n675), .ZN(
        n682) );
  OAI22_X1 U699 ( .A1(n1581), .A2(n79), .B1(n1580), .B2(n76), .ZN(n676) );
  AOI221_X1 U700 ( .B1(n85), .B2(n3995), .C1(n82), .C2(n4029), .A(n676), .ZN(
        n681) );
  OAI22_X1 U701 ( .A1(n1584), .A2(n91), .B1(n1583), .B2(n88), .ZN(n677) );
  AOI221_X1 U702 ( .B1(n97), .B2(n4135), .C1(n94), .C2(n4170), .A(n677), .ZN(
        n680) );
  OAI22_X1 U703 ( .A1(n1587), .A2(n103), .B1(n1586), .B2(n100), .ZN(n678) );
  AOI221_X1 U704 ( .B1(n109), .B2(n4275), .C1(n106), .C2(n4325), .A(n678), 
        .ZN(n679) );
  NAND4_X1 U705 ( .A1(n682), .A2(n681), .A3(n680), .A4(n679), .ZN(n692) );
  OAI22_X1 U706 ( .A1(n1594), .A2(n115), .B1(n1593), .B2(n112), .ZN(n683) );
  AOI221_X1 U707 ( .B1(n121), .B2(n2290), .C1(n118), .C2(n2324), .A(n683), 
        .ZN(n690) );
  OAI22_X1 U708 ( .A1(n1597), .A2(n127), .B1(n1596), .B2(n124), .ZN(n684) );
  AOI221_X1 U709 ( .B1(n133), .B2(n2426), .C1(n130), .C2(n2464), .A(n684), 
        .ZN(n689) );
  OAI22_X1 U710 ( .A1(n1600), .A2(n139), .B1(n1599), .B2(n136), .ZN(n685) );
  AOI221_X1 U711 ( .B1(n145), .B2(n2498), .C1(n142), .C2(n3620), .A(n685), 
        .ZN(n688) );
  OAI22_X1 U712 ( .A1(n1603), .A2(n151), .B1(n1602), .B2(n148), .ZN(n686) );
  AOI221_X1 U713 ( .B1(n157), .B2(n3722), .C1(n154), .C2(n3756), .A(n686), 
        .ZN(n687) );
  NAND4_X1 U714 ( .A1(n690), .A2(n689), .A3(n688), .A4(n687), .ZN(n691) );
  OAI21_X1 U715 ( .B1(n692), .B2(n691), .A(n160), .ZN(n693) );
  OAI21_X1 U716 ( .B1(n163), .B2(n694), .A(n693), .ZN(n2542) );
  OAI22_X1 U717 ( .A1(n1614), .A2(n67), .B1(n1613), .B2(n64), .ZN(n695) );
  AOI221_X1 U718 ( .B1(n73), .B2(n3860), .C1(n70), .C2(n3894), .A(n695), .ZN(
        n702) );
  OAI22_X1 U719 ( .A1(n1617), .A2(n79), .B1(n1616), .B2(n76), .ZN(n696) );
  AOI221_X1 U720 ( .B1(n85), .B2(n3996), .C1(n82), .C2(n4030), .A(n696), .ZN(
        n701) );
  OAI22_X1 U721 ( .A1(n1620), .A2(n91), .B1(n1619), .B2(n88), .ZN(n697) );
  AOI221_X1 U722 ( .B1(n97), .B2(n4136), .C1(n94), .C2(n4171), .A(n697), .ZN(
        n700) );
  OAI22_X1 U723 ( .A1(n1623), .A2(n103), .B1(n1622), .B2(n100), .ZN(n698) );
  AOI221_X1 U724 ( .B1(n109), .B2(n4276), .C1(n106), .C2(n4327), .A(n698), 
        .ZN(n699) );
  NAND4_X1 U725 ( .A1(n702), .A2(n701), .A3(n700), .A4(n699), .ZN(n712) );
  OAI22_X1 U726 ( .A1(n1630), .A2(n115), .B1(n1629), .B2(n112), .ZN(n703) );
  AOI221_X1 U727 ( .B1(n121), .B2(n2291), .C1(n118), .C2(n2325), .A(n703), 
        .ZN(n710) );
  OAI22_X1 U728 ( .A1(n1633), .A2(n127), .B1(n1632), .B2(n124), .ZN(n704) );
  AOI221_X1 U729 ( .B1(n133), .B2(n2427), .C1(n130), .C2(n2465), .A(n704), 
        .ZN(n709) );
  OAI22_X1 U730 ( .A1(n1636), .A2(n139), .B1(n1635), .B2(n136), .ZN(n705) );
  AOI221_X1 U731 ( .B1(n145), .B2(n2499), .C1(n142), .C2(n3621), .A(n705), 
        .ZN(n708) );
  OAI22_X1 U732 ( .A1(n1639), .A2(n151), .B1(n1638), .B2(n148), .ZN(n706) );
  AOI221_X1 U733 ( .B1(n157), .B2(n3723), .C1(n154), .C2(n3757), .A(n706), 
        .ZN(n707) );
  NAND4_X1 U734 ( .A1(n710), .A2(n709), .A3(n708), .A4(n707), .ZN(n711) );
  OAI21_X1 U735 ( .B1(n712), .B2(n711), .A(n160), .ZN(n713) );
  OAI21_X1 U736 ( .B1(n163), .B2(n714), .A(n713), .ZN(n2543) );
  OAI22_X1 U737 ( .A1(n1650), .A2(n67), .B1(n1649), .B2(n64), .ZN(n715) );
  AOI221_X1 U738 ( .B1(n73), .B2(n3861), .C1(n70), .C2(n3895), .A(n715), .ZN(
        n722) );
  OAI22_X1 U739 ( .A1(n1653), .A2(n79), .B1(n1652), .B2(n76), .ZN(n716) );
  AOI221_X1 U740 ( .B1(n85), .B2(n3997), .C1(n82), .C2(n4031), .A(n716), .ZN(
        n721) );
  OAI22_X1 U741 ( .A1(n1656), .A2(n91), .B1(n1655), .B2(n88), .ZN(n717) );
  AOI221_X1 U742 ( .B1(n97), .B2(n4137), .C1(n94), .C2(n4172), .A(n717), .ZN(
        n720) );
  OAI22_X1 U743 ( .A1(n1659), .A2(n103), .B1(n1658), .B2(n100), .ZN(n718) );
  AOI221_X1 U744 ( .B1(n109), .B2(n4277), .C1(n106), .C2(n4329), .A(n718), 
        .ZN(n719) );
  NAND4_X1 U745 ( .A1(n722), .A2(n721), .A3(n720), .A4(n719), .ZN(n732) );
  OAI22_X1 U746 ( .A1(n1666), .A2(n115), .B1(n1665), .B2(n112), .ZN(n723) );
  AOI221_X1 U747 ( .B1(n121), .B2(n2292), .C1(n118), .C2(n2326), .A(n723), 
        .ZN(n730) );
  OAI22_X1 U748 ( .A1(n1669), .A2(n127), .B1(n1668), .B2(n124), .ZN(n724) );
  AOI221_X1 U749 ( .B1(n133), .B2(n2428), .C1(n130), .C2(n2466), .A(n724), 
        .ZN(n729) );
  OAI22_X1 U750 ( .A1(n1672), .A2(n139), .B1(n1671), .B2(n136), .ZN(n725) );
  AOI221_X1 U751 ( .B1(n145), .B2(n2500), .C1(n142), .C2(n3622), .A(n725), 
        .ZN(n728) );
  OAI22_X1 U752 ( .A1(n1675), .A2(n151), .B1(n1674), .B2(n148), .ZN(n726) );
  AOI221_X1 U753 ( .B1(n157), .B2(n3724), .C1(n154), .C2(n3758), .A(n726), 
        .ZN(n727) );
  NAND4_X1 U754 ( .A1(n730), .A2(n729), .A3(n728), .A4(n727), .ZN(n731) );
  OAI21_X1 U755 ( .B1(n732), .B2(n731), .A(n160), .ZN(n733) );
  OAI21_X1 U756 ( .B1(n163), .B2(n734), .A(n733), .ZN(n2544) );
  OAI22_X1 U757 ( .A1(n1686), .A2(n67), .B1(n1685), .B2(n64), .ZN(n735) );
  AOI221_X1 U758 ( .B1(n73), .B2(n3862), .C1(n70), .C2(n3896), .A(n735), .ZN(
        n742) );
  OAI22_X1 U759 ( .A1(n1689), .A2(n79), .B1(n1688), .B2(n76), .ZN(n736) );
  AOI221_X1 U760 ( .B1(n85), .B2(n3998), .C1(n82), .C2(n4032), .A(n736), .ZN(
        n741) );
  OAI22_X1 U761 ( .A1(n1692), .A2(n91), .B1(n1691), .B2(n88), .ZN(n737) );
  AOI221_X1 U762 ( .B1(n97), .B2(n4138), .C1(n94), .C2(n4173), .A(n737), .ZN(
        n740) );
  OAI22_X1 U763 ( .A1(n1695), .A2(n103), .B1(n1694), .B2(n100), .ZN(n738) );
  AOI221_X1 U764 ( .B1(n109), .B2(n4278), .C1(n106), .C2(n4331), .A(n738), 
        .ZN(n739) );
  NAND4_X1 U765 ( .A1(n742), .A2(n741), .A3(n740), .A4(n739), .ZN(n752) );
  OAI22_X1 U766 ( .A1(n1702), .A2(n115), .B1(n1701), .B2(n112), .ZN(n743) );
  AOI221_X1 U767 ( .B1(n121), .B2(n2293), .C1(n118), .C2(n2327), .A(n743), 
        .ZN(n750) );
  OAI22_X1 U768 ( .A1(n1705), .A2(n127), .B1(n1704), .B2(n124), .ZN(n744) );
  AOI221_X1 U769 ( .B1(n133), .B2(n2429), .C1(n130), .C2(n2467), .A(n744), 
        .ZN(n749) );
  OAI22_X1 U770 ( .A1(n1708), .A2(n139), .B1(n1707), .B2(n136), .ZN(n745) );
  AOI221_X1 U771 ( .B1(n145), .B2(n2501), .C1(n142), .C2(n3623), .A(n745), 
        .ZN(n748) );
  OAI22_X1 U772 ( .A1(n1711), .A2(n151), .B1(n1710), .B2(n148), .ZN(n746) );
  AOI221_X1 U773 ( .B1(n157), .B2(n3725), .C1(n154), .C2(n3759), .A(n746), 
        .ZN(n747) );
  NAND4_X1 U774 ( .A1(n750), .A2(n749), .A3(n748), .A4(n747), .ZN(n751) );
  OAI21_X1 U775 ( .B1(n752), .B2(n751), .A(n160), .ZN(n753) );
  OAI21_X1 U776 ( .B1(n163), .B2(n754), .A(n753), .ZN(n2545) );
  OAI22_X1 U777 ( .A1(n1722), .A2(n67), .B1(n1721), .B2(n64), .ZN(n755) );
  AOI221_X1 U778 ( .B1(n73), .B2(n3863), .C1(n70), .C2(n3897), .A(n755), .ZN(
        n762) );
  OAI22_X1 U779 ( .A1(n1725), .A2(n79), .B1(n1724), .B2(n76), .ZN(n756) );
  AOI221_X1 U780 ( .B1(n85), .B2(n3999), .C1(n82), .C2(n4033), .A(n756), .ZN(
        n761) );
  OAI22_X1 U781 ( .A1(n1728), .A2(n91), .B1(n1727), .B2(n88), .ZN(n757) );
  AOI221_X1 U782 ( .B1(n97), .B2(n4139), .C1(n94), .C2(n4174), .A(n757), .ZN(
        n760) );
  OAI22_X1 U783 ( .A1(n1731), .A2(n103), .B1(n1730), .B2(n100), .ZN(n758) );
  AOI221_X1 U784 ( .B1(n109), .B2(n4279), .C1(n106), .C2(n4333), .A(n758), 
        .ZN(n759) );
  NAND4_X1 U785 ( .A1(n762), .A2(n761), .A3(n760), .A4(n759), .ZN(n772) );
  OAI22_X1 U786 ( .A1(n1738), .A2(n115), .B1(n1737), .B2(n112), .ZN(n763) );
  AOI221_X1 U787 ( .B1(n121), .B2(n2294), .C1(n118), .C2(n2328), .A(n763), 
        .ZN(n770) );
  OAI22_X1 U788 ( .A1(n1741), .A2(n127), .B1(n1740), .B2(n124), .ZN(n764) );
  AOI221_X1 U789 ( .B1(n133), .B2(n2430), .C1(n130), .C2(n2468), .A(n764), 
        .ZN(n769) );
  OAI22_X1 U790 ( .A1(n1744), .A2(n139), .B1(n1743), .B2(n136), .ZN(n765) );
  AOI221_X1 U791 ( .B1(n145), .B2(n2502), .C1(n142), .C2(n3624), .A(n765), 
        .ZN(n768) );
  OAI22_X1 U792 ( .A1(n1747), .A2(n151), .B1(n1746), .B2(n148), .ZN(n766) );
  AOI221_X1 U793 ( .B1(n157), .B2(n3726), .C1(n154), .C2(n3760), .A(n766), 
        .ZN(n767) );
  NAND4_X1 U794 ( .A1(n770), .A2(n769), .A3(n768), .A4(n767), .ZN(n771) );
  OAI21_X1 U795 ( .B1(n772), .B2(n771), .A(n160), .ZN(n773) );
  OAI21_X1 U796 ( .B1(n163), .B2(n774), .A(n773), .ZN(n2546) );
  OAI22_X1 U797 ( .A1(n1758), .A2(n67), .B1(n1757), .B2(n64), .ZN(n775) );
  AOI221_X1 U798 ( .B1(n73), .B2(n3864), .C1(n70), .C2(n3898), .A(n775), .ZN(
        n782) );
  OAI22_X1 U799 ( .A1(n1761), .A2(n79), .B1(n1760), .B2(n76), .ZN(n776) );
  AOI221_X1 U800 ( .B1(n85), .B2(n4000), .C1(n82), .C2(n4034), .A(n776), .ZN(
        n781) );
  OAI22_X1 U801 ( .A1(n1764), .A2(n91), .B1(n1763), .B2(n88), .ZN(n777) );
  AOI221_X1 U802 ( .B1(n97), .B2(n4140), .C1(n94), .C2(n4175), .A(n777), .ZN(
        n780) );
  OAI22_X1 U803 ( .A1(n1767), .A2(n103), .B1(n1766), .B2(n100), .ZN(n778) );
  AOI221_X1 U804 ( .B1(n109), .B2(n4280), .C1(n106), .C2(n4335), .A(n778), 
        .ZN(n779) );
  NAND4_X1 U805 ( .A1(n782), .A2(n781), .A3(n780), .A4(n779), .ZN(n792) );
  OAI22_X1 U806 ( .A1(n1774), .A2(n115), .B1(n1773), .B2(n112), .ZN(n783) );
  AOI221_X1 U807 ( .B1(n121), .B2(n2295), .C1(n118), .C2(n2329), .A(n783), 
        .ZN(n790) );
  OAI22_X1 U808 ( .A1(n1777), .A2(n127), .B1(n1776), .B2(n124), .ZN(n784) );
  AOI221_X1 U809 ( .B1(n133), .B2(n2431), .C1(n130), .C2(n2469), .A(n784), 
        .ZN(n789) );
  OAI22_X1 U810 ( .A1(n1780), .A2(n139), .B1(n1779), .B2(n136), .ZN(n785) );
  AOI221_X1 U811 ( .B1(n145), .B2(n2503), .C1(n142), .C2(n3625), .A(n785), 
        .ZN(n788) );
  OAI22_X1 U812 ( .A1(n1783), .A2(n151), .B1(n1782), .B2(n148), .ZN(n786) );
  AOI221_X1 U813 ( .B1(n157), .B2(n3727), .C1(n154), .C2(n3761), .A(n786), 
        .ZN(n787) );
  NAND4_X1 U814 ( .A1(n790), .A2(n789), .A3(n788), .A4(n787), .ZN(n791) );
  OAI21_X1 U815 ( .B1(n792), .B2(n791), .A(n160), .ZN(n793) );
  OAI21_X1 U816 ( .B1(n163), .B2(n794), .A(n793), .ZN(n2547) );
  OAI22_X1 U817 ( .A1(n1794), .A2(n67), .B1(n1793), .B2(n64), .ZN(n795) );
  AOI221_X1 U818 ( .B1(n73), .B2(n3865), .C1(n70), .C2(n3899), .A(n795), .ZN(
        n802) );
  OAI22_X1 U819 ( .A1(n1797), .A2(n79), .B1(n1796), .B2(n76), .ZN(n796) );
  AOI221_X1 U820 ( .B1(n85), .B2(n4001), .C1(n82), .C2(n4035), .A(n796), .ZN(
        n801) );
  OAI22_X1 U821 ( .A1(n1800), .A2(n91), .B1(n1799), .B2(n88), .ZN(n797) );
  AOI221_X1 U822 ( .B1(n97), .B2(n4141), .C1(n94), .C2(n4176), .A(n797), .ZN(
        n800) );
  OAI22_X1 U823 ( .A1(n1803), .A2(n103), .B1(n1802), .B2(n100), .ZN(n798) );
  AOI221_X1 U824 ( .B1(n109), .B2(n4281), .C1(n106), .C2(n4337), .A(n798), 
        .ZN(n799) );
  NAND4_X1 U825 ( .A1(n802), .A2(n801), .A3(n800), .A4(n799), .ZN(n812) );
  OAI22_X1 U826 ( .A1(n1810), .A2(n115), .B1(n1809), .B2(n112), .ZN(n803) );
  AOI221_X1 U827 ( .B1(n121), .B2(n2296), .C1(n118), .C2(n2330), .A(n803), 
        .ZN(n810) );
  OAI22_X1 U828 ( .A1(n1813), .A2(n127), .B1(n1812), .B2(n124), .ZN(n804) );
  AOI221_X1 U829 ( .B1(n133), .B2(n2432), .C1(n130), .C2(n2470), .A(n804), 
        .ZN(n809) );
  OAI22_X1 U830 ( .A1(n1816), .A2(n139), .B1(n1815), .B2(n136), .ZN(n805) );
  AOI221_X1 U831 ( .B1(n145), .B2(n2504), .C1(n142), .C2(n3626), .A(n805), 
        .ZN(n808) );
  OAI22_X1 U832 ( .A1(n1819), .A2(n151), .B1(n1818), .B2(n148), .ZN(n806) );
  AOI221_X1 U833 ( .B1(n157), .B2(n3728), .C1(n154), .C2(n3762), .A(n806), 
        .ZN(n807) );
  NAND4_X1 U834 ( .A1(n810), .A2(n809), .A3(n808), .A4(n807), .ZN(n811) );
  OAI21_X1 U835 ( .B1(n812), .B2(n811), .A(n160), .ZN(n813) );
  OAI21_X1 U836 ( .B1(n163), .B2(n814), .A(n813), .ZN(n2548) );
  OAI22_X1 U837 ( .A1(n1830), .A2(n67), .B1(n1829), .B2(n64), .ZN(n815) );
  AOI221_X1 U838 ( .B1(n73), .B2(n3866), .C1(n70), .C2(n3900), .A(n815), .ZN(
        n822) );
  OAI22_X1 U839 ( .A1(n1833), .A2(n79), .B1(n1832), .B2(n76), .ZN(n816) );
  AOI221_X1 U840 ( .B1(n85), .B2(n4002), .C1(n82), .C2(n4036), .A(n816), .ZN(
        n821) );
  OAI22_X1 U841 ( .A1(n1836), .A2(n91), .B1(n1835), .B2(n88), .ZN(n817) );
  AOI221_X1 U842 ( .B1(n97), .B2(n4142), .C1(n94), .C2(n4177), .A(n817), .ZN(
        n820) );
  OAI22_X1 U843 ( .A1(n1839), .A2(n103), .B1(n1838), .B2(n100), .ZN(n818) );
  AOI221_X1 U844 ( .B1(n109), .B2(n4282), .C1(n106), .C2(n4339), .A(n818), 
        .ZN(n819) );
  NAND4_X1 U845 ( .A1(n822), .A2(n821), .A3(n820), .A4(n819), .ZN(n832) );
  OAI22_X1 U846 ( .A1(n1846), .A2(n115), .B1(n1845), .B2(n112), .ZN(n823) );
  AOI221_X1 U847 ( .B1(n121), .B2(n2297), .C1(n118), .C2(n2331), .A(n823), 
        .ZN(n830) );
  OAI22_X1 U848 ( .A1(n1849), .A2(n127), .B1(n1848), .B2(n124), .ZN(n824) );
  AOI221_X1 U849 ( .B1(n133), .B2(n2433), .C1(n130), .C2(n2471), .A(n824), 
        .ZN(n829) );
  OAI22_X1 U850 ( .A1(n1852), .A2(n139), .B1(n1851), .B2(n136), .ZN(n825) );
  AOI221_X1 U851 ( .B1(n145), .B2(n2505), .C1(n142), .C2(n3627), .A(n825), 
        .ZN(n828) );
  OAI22_X1 U852 ( .A1(n1855), .A2(n151), .B1(n1854), .B2(n148), .ZN(n826) );
  AOI221_X1 U853 ( .B1(n157), .B2(n3729), .C1(n154), .C2(n3763), .A(n826), 
        .ZN(n827) );
  NAND4_X1 U854 ( .A1(n830), .A2(n829), .A3(n828), .A4(n827), .ZN(n831) );
  OAI21_X1 U855 ( .B1(n832), .B2(n831), .A(n160), .ZN(n833) );
  OAI21_X1 U856 ( .B1(n163), .B2(n834), .A(n833), .ZN(n2549) );
  OAI22_X1 U857 ( .A1(n1866), .A2(n67), .B1(n1865), .B2(n64), .ZN(n835) );
  AOI221_X1 U858 ( .B1(n73), .B2(n3867), .C1(n70), .C2(n3901), .A(n835), .ZN(
        n842) );
  OAI22_X1 U859 ( .A1(n1869), .A2(n79), .B1(n1868), .B2(n76), .ZN(n836) );
  AOI221_X1 U860 ( .B1(n85), .B2(n4003), .C1(n82), .C2(n4037), .A(n836), .ZN(
        n841) );
  OAI22_X1 U861 ( .A1(n1872), .A2(n91), .B1(n1871), .B2(n88), .ZN(n837) );
  AOI221_X1 U862 ( .B1(n97), .B2(n4143), .C1(n94), .C2(n4178), .A(n837), .ZN(
        n840) );
  OAI22_X1 U863 ( .A1(n1875), .A2(n103), .B1(n1874), .B2(n100), .ZN(n838) );
  AOI221_X1 U864 ( .B1(n109), .B2(n4283), .C1(n106), .C2(n4341), .A(n838), 
        .ZN(n839) );
  NAND4_X1 U865 ( .A1(n842), .A2(n841), .A3(n840), .A4(n839), .ZN(n852) );
  OAI22_X1 U866 ( .A1(n1882), .A2(n115), .B1(n1881), .B2(n112), .ZN(n843) );
  AOI221_X1 U867 ( .B1(n121), .B2(n2298), .C1(n118), .C2(n2332), .A(n843), 
        .ZN(n850) );
  OAI22_X1 U868 ( .A1(n1885), .A2(n127), .B1(n1884), .B2(n124), .ZN(n844) );
  AOI221_X1 U869 ( .B1(n133), .B2(n2434), .C1(n130), .C2(n2472), .A(n844), 
        .ZN(n849) );
  OAI22_X1 U870 ( .A1(n1888), .A2(n139), .B1(n1887), .B2(n136), .ZN(n845) );
  AOI221_X1 U871 ( .B1(n145), .B2(n2506), .C1(n142), .C2(n3628), .A(n845), 
        .ZN(n848) );
  OAI22_X1 U872 ( .A1(n1891), .A2(n151), .B1(n1890), .B2(n148), .ZN(n846) );
  AOI221_X1 U873 ( .B1(n157), .B2(n3730), .C1(n154), .C2(n3764), .A(n846), 
        .ZN(n847) );
  NAND4_X1 U874 ( .A1(n850), .A2(n849), .A3(n848), .A4(n847), .ZN(n851) );
  OAI21_X1 U875 ( .B1(n852), .B2(n851), .A(n160), .ZN(n853) );
  OAI21_X1 U876 ( .B1(n164), .B2(n854), .A(n853), .ZN(n2550) );
  OAI22_X1 U877 ( .A1(n1902), .A2(n68), .B1(n1901), .B2(n65), .ZN(n855) );
  AOI221_X1 U878 ( .B1(n74), .B2(n3868), .C1(n71), .C2(n3902), .A(n855), .ZN(
        n862) );
  OAI22_X1 U879 ( .A1(n1905), .A2(n80), .B1(n1904), .B2(n77), .ZN(n856) );
  AOI221_X1 U880 ( .B1(n86), .B2(n4004), .C1(n83), .C2(n4038), .A(n856), .ZN(
        n861) );
  OAI22_X1 U881 ( .A1(n1908), .A2(n92), .B1(n1907), .B2(n89), .ZN(n857) );
  AOI221_X1 U882 ( .B1(n98), .B2(n4144), .C1(n95), .C2(n4179), .A(n857), .ZN(
        n860) );
  OAI22_X1 U883 ( .A1(n1911), .A2(n104), .B1(n1910), .B2(n101), .ZN(n858) );
  AOI221_X1 U884 ( .B1(n110), .B2(n4284), .C1(n107), .C2(n4343), .A(n858), 
        .ZN(n859) );
  NAND4_X1 U885 ( .A1(n862), .A2(n861), .A3(n860), .A4(n859), .ZN(n872) );
  OAI22_X1 U886 ( .A1(n1918), .A2(n116), .B1(n1917), .B2(n113), .ZN(n863) );
  AOI221_X1 U887 ( .B1(n122), .B2(n2299), .C1(n119), .C2(n2333), .A(n863), 
        .ZN(n870) );
  OAI22_X1 U888 ( .A1(n1921), .A2(n128), .B1(n1920), .B2(n125), .ZN(n864) );
  AOI221_X1 U889 ( .B1(n134), .B2(n2435), .C1(n131), .C2(n2473), .A(n864), 
        .ZN(n869) );
  OAI22_X1 U890 ( .A1(n1924), .A2(n140), .B1(n1923), .B2(n137), .ZN(n865) );
  AOI221_X1 U891 ( .B1(n146), .B2(n2507), .C1(n143), .C2(n3629), .A(n865), 
        .ZN(n868) );
  OAI22_X1 U892 ( .A1(n1927), .A2(n152), .B1(n1926), .B2(n149), .ZN(n866) );
  AOI221_X1 U893 ( .B1(n158), .B2(n3731), .C1(n155), .C2(n3765), .A(n866), 
        .ZN(n867) );
  NAND4_X1 U894 ( .A1(n870), .A2(n869), .A3(n868), .A4(n867), .ZN(n871) );
  OAI21_X1 U895 ( .B1(n872), .B2(n871), .A(n161), .ZN(n873) );
  OAI21_X1 U896 ( .B1(n164), .B2(n874), .A(n873), .ZN(n2551) );
  OAI22_X1 U897 ( .A1(n1938), .A2(n68), .B1(n1937), .B2(n65), .ZN(n875) );
  AOI221_X1 U898 ( .B1(n74), .B2(n3869), .C1(n71), .C2(n3903), .A(n875), .ZN(
        n882) );
  OAI22_X1 U899 ( .A1(n1941), .A2(n80), .B1(n1940), .B2(n77), .ZN(n876) );
  AOI221_X1 U900 ( .B1(n86), .B2(n4005), .C1(n83), .C2(n4039), .A(n876), .ZN(
        n881) );
  OAI22_X1 U901 ( .A1(n1944), .A2(n92), .B1(n1943), .B2(n89), .ZN(n877) );
  AOI221_X1 U902 ( .B1(n98), .B2(n4145), .C1(n95), .C2(n4180), .A(n877), .ZN(
        n880) );
  OAI22_X1 U903 ( .A1(n1947), .A2(n104), .B1(n1946), .B2(n101), .ZN(n878) );
  AOI221_X1 U904 ( .B1(n110), .B2(n4285), .C1(n107), .C2(n4345), .A(n878), 
        .ZN(n879) );
  NAND4_X1 U905 ( .A1(n882), .A2(n881), .A3(n880), .A4(n879), .ZN(n892) );
  OAI22_X1 U906 ( .A1(n1954), .A2(n116), .B1(n1953), .B2(n113), .ZN(n883) );
  AOI221_X1 U907 ( .B1(n122), .B2(n2300), .C1(n119), .C2(n2334), .A(n883), 
        .ZN(n890) );
  OAI22_X1 U908 ( .A1(n1957), .A2(n128), .B1(n1956), .B2(n125), .ZN(n884) );
  AOI221_X1 U909 ( .B1(n134), .B2(n2436), .C1(n131), .C2(n2474), .A(n884), 
        .ZN(n889) );
  OAI22_X1 U910 ( .A1(n1960), .A2(n140), .B1(n1959), .B2(n137), .ZN(n885) );
  AOI221_X1 U911 ( .B1(n146), .B2(n2508), .C1(n143), .C2(n3630), .A(n885), 
        .ZN(n888) );
  OAI22_X1 U912 ( .A1(n1963), .A2(n152), .B1(n1962), .B2(n149), .ZN(n886) );
  AOI221_X1 U913 ( .B1(n158), .B2(n3732), .C1(n155), .C2(n3766), .A(n886), 
        .ZN(n887) );
  NAND4_X1 U914 ( .A1(n890), .A2(n889), .A3(n888), .A4(n887), .ZN(n891) );
  OAI21_X1 U915 ( .B1(n892), .B2(n891), .A(n161), .ZN(n893) );
  OAI21_X1 U916 ( .B1(n164), .B2(n894), .A(n893), .ZN(n2552) );
  OAI22_X1 U917 ( .A1(n1974), .A2(n68), .B1(n1973), .B2(n65), .ZN(n895) );
  AOI221_X1 U918 ( .B1(n74), .B2(n3870), .C1(n71), .C2(n3904), .A(n895), .ZN(
        n902) );
  OAI22_X1 U919 ( .A1(n1977), .A2(n80), .B1(n1976), .B2(n77), .ZN(n896) );
  AOI221_X1 U920 ( .B1(n86), .B2(n4006), .C1(n83), .C2(n4040), .A(n896), .ZN(
        n901) );
  OAI22_X1 U921 ( .A1(n1980), .A2(n92), .B1(n1979), .B2(n89), .ZN(n897) );
  AOI221_X1 U922 ( .B1(n98), .B2(n4146), .C1(n95), .C2(n4181), .A(n897), .ZN(
        n900) );
  OAI22_X1 U923 ( .A1(n1983), .A2(n104), .B1(n1982), .B2(n101), .ZN(n898) );
  AOI221_X1 U924 ( .B1(n110), .B2(n4286), .C1(n107), .C2(n4347), .A(n898), 
        .ZN(n899) );
  NAND4_X1 U925 ( .A1(n902), .A2(n901), .A3(n900), .A4(n899), .ZN(n912) );
  OAI22_X1 U926 ( .A1(n1990), .A2(n116), .B1(n1989), .B2(n113), .ZN(n903) );
  AOI221_X1 U927 ( .B1(n122), .B2(n2301), .C1(n119), .C2(n2335), .A(n903), 
        .ZN(n910) );
  OAI22_X1 U928 ( .A1(n1993), .A2(n128), .B1(n1992), .B2(n125), .ZN(n904) );
  AOI221_X1 U929 ( .B1(n134), .B2(n2437), .C1(n131), .C2(n2475), .A(n904), 
        .ZN(n909) );
  OAI22_X1 U930 ( .A1(n1996), .A2(n140), .B1(n1995), .B2(n137), .ZN(n905) );
  AOI221_X1 U931 ( .B1(n146), .B2(n2509), .C1(n143), .C2(n3631), .A(n905), 
        .ZN(n908) );
  OAI22_X1 U932 ( .A1(n1999), .A2(n152), .B1(n1998), .B2(n149), .ZN(n906) );
  AOI221_X1 U933 ( .B1(n158), .B2(n3733), .C1(n155), .C2(n3767), .A(n906), 
        .ZN(n907) );
  NAND4_X1 U934 ( .A1(n910), .A2(n909), .A3(n908), .A4(n907), .ZN(n911) );
  OAI21_X1 U935 ( .B1(n912), .B2(n911), .A(n161), .ZN(n913) );
  OAI21_X1 U936 ( .B1(n164), .B2(n914), .A(n913), .ZN(n2553) );
  OAI22_X1 U937 ( .A1(n2010), .A2(n68), .B1(n2009), .B2(n65), .ZN(n915) );
  AOI221_X1 U938 ( .B1(n74), .B2(n3871), .C1(n71), .C2(n3905), .A(n915), .ZN(
        n922) );
  OAI22_X1 U939 ( .A1(n2013), .A2(n80), .B1(n2012), .B2(n77), .ZN(n916) );
  AOI221_X1 U940 ( .B1(n86), .B2(n4007), .C1(n83), .C2(n4041), .A(n916), .ZN(
        n921) );
  OAI22_X1 U941 ( .A1(n2016), .A2(n92), .B1(n2015), .B2(n89), .ZN(n917) );
  AOI221_X1 U942 ( .B1(n98), .B2(n4147), .C1(n95), .C2(n4182), .A(n917), .ZN(
        n920) );
  OAI22_X1 U943 ( .A1(n2019), .A2(n104), .B1(n2018), .B2(n101), .ZN(n918) );
  AOI221_X1 U944 ( .B1(n110), .B2(n4287), .C1(n107), .C2(n4349), .A(n918), 
        .ZN(n919) );
  NAND4_X1 U945 ( .A1(n922), .A2(n921), .A3(n920), .A4(n919), .ZN(n932) );
  OAI22_X1 U946 ( .A1(n2026), .A2(n116), .B1(n2025), .B2(n113), .ZN(n923) );
  AOI221_X1 U947 ( .B1(n122), .B2(n2302), .C1(n119), .C2(n2336), .A(n923), 
        .ZN(n930) );
  OAI22_X1 U948 ( .A1(n2029), .A2(n128), .B1(n2028), .B2(n125), .ZN(n924) );
  AOI221_X1 U949 ( .B1(n134), .B2(n2438), .C1(n131), .C2(n2476), .A(n924), 
        .ZN(n929) );
  OAI22_X1 U950 ( .A1(n2032), .A2(n140), .B1(n2031), .B2(n137), .ZN(n925) );
  AOI221_X1 U951 ( .B1(n146), .B2(n2510), .C1(n143), .C2(n3632), .A(n925), 
        .ZN(n928) );
  OAI22_X1 U952 ( .A1(n2035), .A2(n152), .B1(n2034), .B2(n149), .ZN(n926) );
  AOI221_X1 U953 ( .B1(n158), .B2(n3734), .C1(n155), .C2(n3768), .A(n926), 
        .ZN(n927) );
  NAND4_X1 U954 ( .A1(n930), .A2(n929), .A3(n928), .A4(n927), .ZN(n931) );
  OAI21_X1 U955 ( .B1(n932), .B2(n931), .A(n161), .ZN(n933) );
  OAI21_X1 U956 ( .B1(n164), .B2(n934), .A(n933), .ZN(n2554) );
  OAI22_X1 U957 ( .A1(n2046), .A2(n68), .B1(n2045), .B2(n65), .ZN(n935) );
  AOI221_X1 U958 ( .B1(n74), .B2(n3872), .C1(n71), .C2(n3906), .A(n935), .ZN(
        n942) );
  OAI22_X1 U959 ( .A1(n2049), .A2(n80), .B1(n2048), .B2(n77), .ZN(n936) );
  AOI221_X1 U960 ( .B1(n86), .B2(n4008), .C1(n83), .C2(n4042), .A(n936), .ZN(
        n941) );
  OAI22_X1 U961 ( .A1(n2052), .A2(n92), .B1(n2051), .B2(n89), .ZN(n937) );
  AOI221_X1 U962 ( .B1(n98), .B2(n4148), .C1(n95), .C2(n4183), .A(n937), .ZN(
        n940) );
  OAI22_X1 U963 ( .A1(n2055), .A2(n104), .B1(n2054), .B2(n101), .ZN(n938) );
  AOI221_X1 U964 ( .B1(n110), .B2(n4288), .C1(n107), .C2(n4351), .A(n938), 
        .ZN(n939) );
  NAND4_X1 U965 ( .A1(n942), .A2(n941), .A3(n940), .A4(n939), .ZN(n952) );
  OAI22_X1 U966 ( .A1(n2062), .A2(n116), .B1(n2061), .B2(n113), .ZN(n943) );
  AOI221_X1 U967 ( .B1(n122), .B2(n2303), .C1(n119), .C2(n2337), .A(n943), 
        .ZN(n950) );
  OAI22_X1 U968 ( .A1(n2065), .A2(n128), .B1(n2064), .B2(n125), .ZN(n944) );
  AOI221_X1 U969 ( .B1(n134), .B2(n2439), .C1(n131), .C2(n2477), .A(n944), 
        .ZN(n949) );
  OAI22_X1 U970 ( .A1(n2068), .A2(n140), .B1(n2067), .B2(n137), .ZN(n945) );
  AOI221_X1 U971 ( .B1(n146), .B2(n2511), .C1(n143), .C2(n3633), .A(n945), 
        .ZN(n948) );
  OAI22_X1 U972 ( .A1(n2071), .A2(n152), .B1(n2070), .B2(n149), .ZN(n946) );
  AOI221_X1 U973 ( .B1(n158), .B2(n3735), .C1(n155), .C2(n3769), .A(n946), 
        .ZN(n947) );
  NAND4_X1 U974 ( .A1(n950), .A2(n949), .A3(n948), .A4(n947), .ZN(n951) );
  OAI21_X1 U975 ( .B1(n952), .B2(n951), .A(n161), .ZN(n953) );
  OAI21_X1 U976 ( .B1(n164), .B2(n954), .A(n953), .ZN(n2555) );
  OAI22_X1 U977 ( .A1(n2082), .A2(n68), .B1(n2081), .B2(n65), .ZN(n955) );
  AOI221_X1 U978 ( .B1(n74), .B2(n3873), .C1(n71), .C2(n3907), .A(n955), .ZN(
        n962) );
  OAI22_X1 U979 ( .A1(n2085), .A2(n80), .B1(n2084), .B2(n77), .ZN(n956) );
  AOI221_X1 U980 ( .B1(n86), .B2(n4009), .C1(n83), .C2(n4043), .A(n956), .ZN(
        n961) );
  OAI22_X1 U981 ( .A1(n2088), .A2(n92), .B1(n2087), .B2(n89), .ZN(n957) );
  AOI221_X1 U982 ( .B1(n98), .B2(n4149), .C1(n95), .C2(n4184), .A(n957), .ZN(
        n960) );
  OAI22_X1 U983 ( .A1(n2091), .A2(n104), .B1(n2090), .B2(n101), .ZN(n958) );
  AOI221_X1 U984 ( .B1(n110), .B2(n4289), .C1(n107), .C2(n4353), .A(n958), 
        .ZN(n959) );
  NAND4_X1 U985 ( .A1(n962), .A2(n961), .A3(n960), .A4(n959), .ZN(n972) );
  OAI22_X1 U986 ( .A1(n2098), .A2(n116), .B1(n2097), .B2(n113), .ZN(n963) );
  AOI221_X1 U987 ( .B1(n122), .B2(n2304), .C1(n119), .C2(n2338), .A(n963), 
        .ZN(n970) );
  OAI22_X1 U988 ( .A1(n2101), .A2(n128), .B1(n2100), .B2(n125), .ZN(n964) );
  AOI221_X1 U989 ( .B1(n134), .B2(n2440), .C1(n131), .C2(n2478), .A(n964), 
        .ZN(n969) );
  OAI22_X1 U990 ( .A1(n2104), .A2(n140), .B1(n2103), .B2(n137), .ZN(n965) );
  AOI221_X1 U991 ( .B1(n146), .B2(n2512), .C1(n143), .C2(n3634), .A(n965), 
        .ZN(n968) );
  OAI22_X1 U992 ( .A1(n2107), .A2(n152), .B1(n2106), .B2(n149), .ZN(n966) );
  AOI221_X1 U993 ( .B1(n158), .B2(n3736), .C1(n155), .C2(n3770), .A(n966), 
        .ZN(n967) );
  NAND4_X1 U994 ( .A1(n970), .A2(n969), .A3(n968), .A4(n967), .ZN(n971) );
  OAI21_X1 U995 ( .B1(n972), .B2(n971), .A(n161), .ZN(n973) );
  OAI21_X1 U996 ( .B1(n164), .B2(n974), .A(n973), .ZN(n2556) );
  OAI22_X1 U997 ( .A1(n2118), .A2(n68), .B1(n2117), .B2(n65), .ZN(n975) );
  AOI221_X1 U998 ( .B1(n74), .B2(n3874), .C1(n71), .C2(n3908), .A(n975), .ZN(
        n982) );
  OAI22_X1 U999 ( .A1(n2121), .A2(n80), .B1(n2120), .B2(n77), .ZN(n976) );
  AOI221_X1 U1000 ( .B1(n86), .B2(n4010), .C1(n83), .C2(n4044), .A(n976), .ZN(
        n981) );
  OAI22_X1 U1001 ( .A1(n2124), .A2(n92), .B1(n2123), .B2(n89), .ZN(n977) );
  AOI221_X1 U1002 ( .B1(n98), .B2(n4150), .C1(n95), .C2(n4185), .A(n977), .ZN(
        n980) );
  OAI22_X1 U1003 ( .A1(n2127), .A2(n104), .B1(n2126), .B2(n101), .ZN(n978) );
  AOI221_X1 U1004 ( .B1(n110), .B2(n4290), .C1(n107), .C2(n4355), .A(n978), 
        .ZN(n979) );
  NAND4_X1 U1005 ( .A1(n982), .A2(n981), .A3(n980), .A4(n979), .ZN(n992) );
  OAI22_X1 U1006 ( .A1(n2134), .A2(n116), .B1(n2133), .B2(n113), .ZN(n983) );
  AOI221_X1 U1007 ( .B1(n122), .B2(n2305), .C1(n119), .C2(n2339), .A(n983), 
        .ZN(n990) );
  OAI22_X1 U1008 ( .A1(n2137), .A2(n128), .B1(n2136), .B2(n125), .ZN(n984) );
  AOI221_X1 U1009 ( .B1(n134), .B2(n2441), .C1(n131), .C2(n2479), .A(n984), 
        .ZN(n989) );
  OAI22_X1 U1010 ( .A1(n2140), .A2(n140), .B1(n2139), .B2(n137), .ZN(n985) );
  AOI221_X1 U1011 ( .B1(n146), .B2(n2513), .C1(n143), .C2(n3635), .A(n985), 
        .ZN(n988) );
  OAI22_X1 U1012 ( .A1(n2143), .A2(n152), .B1(n2142), .B2(n149), .ZN(n986) );
  AOI221_X1 U1013 ( .B1(n158), .B2(n3737), .C1(n155), .C2(n3771), .A(n986), 
        .ZN(n987) );
  NAND4_X1 U1014 ( .A1(n990), .A2(n989), .A3(n988), .A4(n987), .ZN(n991) );
  OAI21_X1 U1015 ( .B1(n992), .B2(n991), .A(n161), .ZN(n993) );
  OAI21_X1 U1016 ( .B1(n164), .B2(n994), .A(n993), .ZN(n2557) );
  OAI22_X1 U1017 ( .A1(n2155), .A2(n68), .B1(n2153), .B2(n65), .ZN(n997) );
  AOI221_X1 U1018 ( .B1(n74), .B2(n3876), .C1(n71), .C2(n3910), .A(n997), .ZN(
        n1010) );
  OAI22_X1 U1019 ( .A1(n2160), .A2(n80), .B1(n2158), .B2(n77), .ZN(n1000) );
  AOI221_X1 U1020 ( .B1(n86), .B2(n4012), .C1(n83), .C2(n4046), .A(n1000), 
        .ZN(n1009) );
  OAI22_X1 U1021 ( .A1(n2165), .A2(n92), .B1(n2163), .B2(n89), .ZN(n1003) );
  AOI221_X1 U1022 ( .B1(n98), .B2(n4152), .C1(n95), .C2(n4187), .A(n1003), 
        .ZN(n1008) );
  OAI22_X1 U1023 ( .A1(n2170), .A2(n104), .B1(n2168), .B2(n101), .ZN(n1006) );
  AOI221_X1 U1024 ( .B1(n110), .B2(n4292), .C1(n107), .C2(n4358), .A(n1006), 
        .ZN(n1007) );
  NAND4_X1 U1025 ( .A1(n1010), .A2(n1009), .A3(n1008), .A4(n1007), .ZN(n1028)
         );
  OAI22_X1 U1026 ( .A1(n2179), .A2(n116), .B1(n2177), .B2(n113), .ZN(n1013) );
  AOI221_X1 U1027 ( .B1(n122), .B2(n2307), .C1(n119), .C2(n2341), .A(n1013), 
        .ZN(n1026) );
  OAI22_X1 U1028 ( .A1(n2184), .A2(n128), .B1(n2182), .B2(n125), .ZN(n1016) );
  AOI221_X1 U1029 ( .B1(n134), .B2(n2443), .C1(n131), .C2(n2481), .A(n1016), 
        .ZN(n1025) );
  OAI22_X1 U1030 ( .A1(n2189), .A2(n140), .B1(n2187), .B2(n137), .ZN(n1019) );
  AOI221_X1 U1031 ( .B1(n146), .B2(n2515), .C1(n143), .C2(n3637), .A(n1019), 
        .ZN(n1024) );
  OAI22_X1 U1032 ( .A1(n2194), .A2(n152), .B1(n2192), .B2(n149), .ZN(n1022) );
  AOI221_X1 U1033 ( .B1(n158), .B2(n3739), .C1(n155), .C2(n3773), .A(n1022), 
        .ZN(n1023) );
  NAND4_X1 U1034 ( .A1(n1026), .A2(n1025), .A3(n1024), .A4(n1023), .ZN(n1027)
         );
  OAI21_X1 U1035 ( .B1(n1028), .B2(n1027), .A(n161), .ZN(n1029) );
  OAI21_X1 U1036 ( .B1(n164), .B2(n1030), .A(n1029), .ZN(n2558) );
  OR2_X1 U1037 ( .A1(RD1), .A2(n369), .ZN(n2205) );
  INV_X1 U1038 ( .A(ADD_RD1[4]), .ZN(n1040) );
  INV_X1 U1039 ( .A(ADD_RD1[0]), .ZN(n1058) );
  INV_X1 U1040 ( .A(ADD_RD1[1]), .ZN(n1036) );
  NAND2_X1 U1041 ( .A1(n58), .A2(n47), .ZN(n2156) );
  NAND2_X1 U1042 ( .A1(n59), .A2(n47), .ZN(n2154) );
  OAI22_X1 U1043 ( .A1(n168), .A2(n1033), .B1(n165), .B2(n1032), .ZN(n1034) );
  AOI221_X1 U1044 ( .B1(n174), .B2(n3844), .C1(n171), .C2(n3878), .A(n1034), 
        .ZN(n1050) );
  INV_X1 U1045 ( .A(ADD_RD1[2]), .ZN(n1035) );
  NAND2_X1 U1046 ( .A1(n58), .A2(n10), .ZN(n2161) );
  NAND2_X1 U1047 ( .A1(n59), .A2(n10), .ZN(n2159) );
  OAI22_X1 U1048 ( .A1(n180), .A2(n1038), .B1(n177), .B2(n1037), .ZN(n1039) );
  AOI221_X1 U1049 ( .B1(n186), .B2(n3980), .C1(n183), .C2(n4014), .A(n1039), 
        .ZN(n1049) );
  INV_X1 U1050 ( .A(ADD_RD1[3]), .ZN(n1057) );
  NAND2_X1 U1051 ( .A1(n57), .A2(n47), .ZN(n2166) );
  NAND2_X1 U1052 ( .A1(n14), .A2(n47), .ZN(n2164) );
  OAI22_X1 U1053 ( .A1(n192), .A2(n1042), .B1(n189), .B2(n1041), .ZN(n1043) );
  AOI221_X1 U1054 ( .B1(n198), .B2(n4120), .C1(n195), .C2(n4155), .A(n1043), 
        .ZN(n1048) );
  NAND2_X1 U1055 ( .A1(n57), .A2(n10), .ZN(n2171) );
  NAND2_X1 U1056 ( .A1(n14), .A2(n10), .ZN(n2169) );
  OAI22_X1 U1057 ( .A1(n204), .A2(n1045), .B1(n201), .B2(n1044), .ZN(n1046) );
  AOI221_X1 U1058 ( .B1(n210), .B2(n4260), .C1(n207), .C2(n4295), .A(n1046), 
        .ZN(n1047) );
  NAND4_X1 U1059 ( .A1(n1050), .A2(n1049), .A3(n1048), .A4(n1047), .ZN(n1070)
         );
  NAND2_X1 U1060 ( .A1(n3), .A2(n49), .ZN(n2180) );
  NAND2_X1 U1061 ( .A1(n3), .A2(n12), .ZN(n2178) );
  OAI22_X1 U1062 ( .A1(n216), .A2(n1052), .B1(n213), .B2(n1051), .ZN(n1053) );
  AOI221_X1 U1063 ( .B1(n222), .B2(n2275), .C1(n219), .C2(n2309), .A(n1053), 
        .ZN(n1068) );
  NAND2_X1 U1064 ( .A1(n4), .A2(n49), .ZN(n2185) );
  NAND2_X1 U1065 ( .A1(n4), .A2(n12), .ZN(n2183) );
  OAI22_X1 U1066 ( .A1(n228), .A2(n1055), .B1(n225), .B2(n1054), .ZN(n1056) );
  AOI221_X1 U1067 ( .B1(n234), .B2(n2411), .C1(n231), .C2(n2449), .A(n1056), 
        .ZN(n1067) );
  NAND2_X1 U1068 ( .A1(n56), .A2(n47), .ZN(n2190) );
  NAND2_X1 U1069 ( .A1(n55), .A2(n47), .ZN(n2188) );
  OAI22_X1 U1070 ( .A1(n240), .A2(n1060), .B1(n237), .B2(n1059), .ZN(n1061) );
  AOI221_X1 U1071 ( .B1(n246), .B2(n2483), .C1(n243), .C2(n2517), .A(n1061), 
        .ZN(n1066) );
  NAND2_X1 U1072 ( .A1(n56), .A2(n10), .ZN(n2195) );
  NAND2_X1 U1073 ( .A1(n55), .A2(n10), .ZN(n2193) );
  OAI22_X1 U1074 ( .A1(n252), .A2(n1063), .B1(n249), .B2(n1062), .ZN(n1064) );
  AOI221_X1 U1075 ( .B1(n258), .B2(n3707), .C1(n255), .C2(n3741), .A(n1064), 
        .ZN(n1065) );
  NAND4_X1 U1076 ( .A1(n1068), .A2(n1067), .A3(n1066), .A4(n1065), .ZN(n1069)
         );
  OAI21_X1 U1077 ( .B1(n1070), .B2(n1069), .A(n261), .ZN(n1071) );
  OAI21_X1 U1078 ( .B1(n264), .B2(n1072), .A(n1071), .ZN(n2559) );
  OAI22_X1 U1079 ( .A1(n168), .A2(n1074), .B1(n165), .B2(n1073), .ZN(n1075) );
  AOI221_X1 U1080 ( .B1(n174), .B2(n3845), .C1(n171), .C2(n3879), .A(n1075), 
        .ZN(n1088) );
  OAI22_X1 U1081 ( .A1(n180), .A2(n1077), .B1(n177), .B2(n1076), .ZN(n1078) );
  AOI221_X1 U1082 ( .B1(n186), .B2(n3981), .C1(n183), .C2(n4015), .A(n1078), 
        .ZN(n1087) );
  OAI22_X1 U1083 ( .A1(n192), .A2(n1080), .B1(n189), .B2(n1079), .ZN(n1081) );
  AOI221_X1 U1084 ( .B1(n198), .B2(n4121), .C1(n195), .C2(n4156), .A(n1081), 
        .ZN(n1086) );
  OAI22_X1 U1085 ( .A1(n204), .A2(n1083), .B1(n201), .B2(n1082), .ZN(n1084) );
  AOI221_X1 U1086 ( .B1(n210), .B2(n4261), .C1(n207), .C2(n4297), .A(n1084), 
        .ZN(n1085) );
  NAND4_X1 U1087 ( .A1(n1088), .A2(n1087), .A3(n1086), .A4(n1085), .ZN(n1106)
         );
  OAI22_X1 U1088 ( .A1(n216), .A2(n1090), .B1(n213), .B2(n1089), .ZN(n1091) );
  AOI221_X1 U1089 ( .B1(n222), .B2(n2276), .C1(n219), .C2(n2310), .A(n1091), 
        .ZN(n1104) );
  OAI22_X1 U1090 ( .A1(n228), .A2(n1093), .B1(n225), .B2(n1092), .ZN(n1094) );
  AOI221_X1 U1091 ( .B1(n234), .B2(n2412), .C1(n231), .C2(n2450), .A(n1094), 
        .ZN(n1103) );
  OAI22_X1 U1092 ( .A1(n240), .A2(n1096), .B1(n237), .B2(n1095), .ZN(n1097) );
  AOI221_X1 U1093 ( .B1(n246), .B2(n2484), .C1(n243), .C2(n2518), .A(n1097), 
        .ZN(n1102) );
  OAI22_X1 U1094 ( .A1(n252), .A2(n1099), .B1(n249), .B2(n1098), .ZN(n1100) );
  AOI221_X1 U1095 ( .B1(n258), .B2(n3708), .C1(n255), .C2(n3742), .A(n1100), 
        .ZN(n1101) );
  NAND4_X1 U1096 ( .A1(n1104), .A2(n1103), .A3(n1102), .A4(n1101), .ZN(n1105)
         );
  OAI21_X1 U1097 ( .B1(n1106), .B2(n1105), .A(n261), .ZN(n1107) );
  OAI21_X1 U1098 ( .B1(n264), .B2(n1108), .A(n1107), .ZN(n2560) );
  OAI22_X1 U1099 ( .A1(n168), .A2(n1110), .B1(n165), .B2(n1109), .ZN(n1111) );
  AOI221_X1 U1100 ( .B1(n174), .B2(n3846), .C1(n171), .C2(n3880), .A(n1111), 
        .ZN(n1124) );
  OAI22_X1 U1101 ( .A1(n180), .A2(n1113), .B1(n177), .B2(n1112), .ZN(n1114) );
  AOI221_X1 U1102 ( .B1(n186), .B2(n3982), .C1(n183), .C2(n4016), .A(n1114), 
        .ZN(n1123) );
  OAI22_X1 U1103 ( .A1(n192), .A2(n1116), .B1(n189), .B2(n1115), .ZN(n1117) );
  AOI221_X1 U1104 ( .B1(n198), .B2(n4122), .C1(n195), .C2(n4157), .A(n1117), 
        .ZN(n1122) );
  OAI22_X1 U1105 ( .A1(n204), .A2(n1119), .B1(n201), .B2(n1118), .ZN(n1120) );
  AOI221_X1 U1106 ( .B1(n210), .B2(n4262), .C1(n207), .C2(n4299), .A(n1120), 
        .ZN(n1121) );
  NAND4_X1 U1107 ( .A1(n1124), .A2(n1123), .A3(n1122), .A4(n1121), .ZN(n1142)
         );
  OAI22_X1 U1108 ( .A1(n216), .A2(n1126), .B1(n213), .B2(n1125), .ZN(n1127) );
  AOI221_X1 U1109 ( .B1(n222), .B2(n2277), .C1(n219), .C2(n2311), .A(n1127), 
        .ZN(n1140) );
  OAI22_X1 U1110 ( .A1(n228), .A2(n1129), .B1(n225), .B2(n1128), .ZN(n1130) );
  AOI221_X1 U1111 ( .B1(n234), .B2(n2413), .C1(n231), .C2(n2451), .A(n1130), 
        .ZN(n1139) );
  OAI22_X1 U1112 ( .A1(n240), .A2(n1132), .B1(n237), .B2(n1131), .ZN(n1133) );
  AOI221_X1 U1113 ( .B1(n246), .B2(n2485), .C1(n243), .C2(n2519), .A(n1133), 
        .ZN(n1138) );
  OAI22_X1 U1114 ( .A1(n252), .A2(n1135), .B1(n249), .B2(n1134), .ZN(n1136) );
  AOI221_X1 U1115 ( .B1(n258), .B2(n3709), .C1(n255), .C2(n3743), .A(n1136), 
        .ZN(n1137) );
  NAND4_X1 U1116 ( .A1(n1140), .A2(n1139), .A3(n1138), .A4(n1137), .ZN(n1141)
         );
  OAI21_X1 U1117 ( .B1(n1142), .B2(n1141), .A(n261), .ZN(n1143) );
  OAI21_X1 U1118 ( .B1(n264), .B2(n1144), .A(n1143), .ZN(n2561) );
  OAI22_X1 U1119 ( .A1(n168), .A2(n1146), .B1(n165), .B2(n1145), .ZN(n1147) );
  AOI221_X1 U1120 ( .B1(n174), .B2(n3847), .C1(n171), .C2(n3881), .A(n1147), 
        .ZN(n1160) );
  OAI22_X1 U1121 ( .A1(n180), .A2(n1149), .B1(n177), .B2(n1148), .ZN(n1150) );
  AOI221_X1 U1122 ( .B1(n186), .B2(n3983), .C1(n183), .C2(n4017), .A(n1150), 
        .ZN(n1159) );
  OAI22_X1 U1123 ( .A1(n192), .A2(n1152), .B1(n189), .B2(n1151), .ZN(n1153) );
  AOI221_X1 U1124 ( .B1(n198), .B2(n4123), .C1(n195), .C2(n4158), .A(n1153), 
        .ZN(n1158) );
  OAI22_X1 U1125 ( .A1(n204), .A2(n1155), .B1(n201), .B2(n1154), .ZN(n1156) );
  AOI221_X1 U1126 ( .B1(n210), .B2(n4263), .C1(n207), .C2(n4301), .A(n1156), 
        .ZN(n1157) );
  NAND4_X1 U1127 ( .A1(n1160), .A2(n1159), .A3(n1158), .A4(n1157), .ZN(n1178)
         );
  OAI22_X1 U1128 ( .A1(n216), .A2(n1162), .B1(n213), .B2(n1161), .ZN(n1163) );
  AOI221_X1 U1129 ( .B1(n222), .B2(n2278), .C1(n219), .C2(n2312), .A(n1163), 
        .ZN(n1176) );
  OAI22_X1 U1130 ( .A1(n228), .A2(n1165), .B1(n225), .B2(n1164), .ZN(n1166) );
  AOI221_X1 U1131 ( .B1(n234), .B2(n2414), .C1(n231), .C2(n2452), .A(n1166), 
        .ZN(n1175) );
  OAI22_X1 U1132 ( .A1(n240), .A2(n1168), .B1(n237), .B2(n1167), .ZN(n1169) );
  AOI221_X1 U1133 ( .B1(n246), .B2(n2486), .C1(n243), .C2(n2520), .A(n1169), 
        .ZN(n1174) );
  OAI22_X1 U1134 ( .A1(n252), .A2(n1171), .B1(n249), .B2(n1170), .ZN(n1172) );
  AOI221_X1 U1135 ( .B1(n258), .B2(n3710), .C1(n255), .C2(n3744), .A(n1172), 
        .ZN(n1173) );
  NAND4_X1 U1136 ( .A1(n1176), .A2(n1175), .A3(n1174), .A4(n1173), .ZN(n1177)
         );
  OAI21_X1 U1137 ( .B1(n1178), .B2(n1177), .A(n261), .ZN(n1179) );
  OAI21_X1 U1138 ( .B1(n264), .B2(n1180), .A(n1179), .ZN(n2562) );
  OAI22_X1 U1139 ( .A1(n168), .A2(n1182), .B1(n165), .B2(n1181), .ZN(n1183) );
  AOI221_X1 U1140 ( .B1(n174), .B2(n3848), .C1(n171), .C2(n3882), .A(n1183), 
        .ZN(n1196) );
  OAI22_X1 U1141 ( .A1(n180), .A2(n1185), .B1(n177), .B2(n1184), .ZN(n1186) );
  AOI221_X1 U1142 ( .B1(n186), .B2(n3984), .C1(n183), .C2(n4018), .A(n1186), 
        .ZN(n1195) );
  OAI22_X1 U1143 ( .A1(n192), .A2(n1188), .B1(n189), .B2(n1187), .ZN(n1189) );
  AOI221_X1 U1144 ( .B1(n198), .B2(n4124), .C1(n195), .C2(n4159), .A(n1189), 
        .ZN(n1194) );
  OAI22_X1 U1145 ( .A1(n204), .A2(n1191), .B1(n201), .B2(n1190), .ZN(n1192) );
  AOI221_X1 U1146 ( .B1(n210), .B2(n4264), .C1(n207), .C2(n4303), .A(n1192), 
        .ZN(n1193) );
  NAND4_X1 U1147 ( .A1(n1196), .A2(n1195), .A3(n1194), .A4(n1193), .ZN(n1214)
         );
  OAI22_X1 U1148 ( .A1(n216), .A2(n1198), .B1(n213), .B2(n1197), .ZN(n1199) );
  AOI221_X1 U1149 ( .B1(n222), .B2(n2279), .C1(n219), .C2(n2313), .A(n1199), 
        .ZN(n1212) );
  OAI22_X1 U1150 ( .A1(n228), .A2(n1201), .B1(n225), .B2(n1200), .ZN(n1202) );
  AOI221_X1 U1151 ( .B1(n234), .B2(n2415), .C1(n231), .C2(n2453), .A(n1202), 
        .ZN(n1211) );
  OAI22_X1 U1152 ( .A1(n240), .A2(n1204), .B1(n237), .B2(n1203), .ZN(n1205) );
  AOI221_X1 U1153 ( .B1(n246), .B2(n2487), .C1(n243), .C2(n2521), .A(n1205), 
        .ZN(n1210) );
  OAI22_X1 U1154 ( .A1(n252), .A2(n1207), .B1(n249), .B2(n1206), .ZN(n1208) );
  AOI221_X1 U1155 ( .B1(n258), .B2(n3711), .C1(n255), .C2(n3745), .A(n1208), 
        .ZN(n1209) );
  NAND4_X1 U1156 ( .A1(n1212), .A2(n1211), .A3(n1210), .A4(n1209), .ZN(n1213)
         );
  OAI21_X1 U1157 ( .B1(n1214), .B2(n1213), .A(n261), .ZN(n1215) );
  OAI21_X1 U1158 ( .B1(n264), .B2(n1216), .A(n1215), .ZN(n2563) );
  OAI22_X1 U1159 ( .A1(n168), .A2(n1218), .B1(n165), .B2(n1217), .ZN(n1219) );
  AOI221_X1 U1160 ( .B1(n174), .B2(n3849), .C1(n171), .C2(n3883), .A(n1219), 
        .ZN(n1232) );
  OAI22_X1 U1161 ( .A1(n180), .A2(n1221), .B1(n177), .B2(n1220), .ZN(n1222) );
  AOI221_X1 U1162 ( .B1(n186), .B2(n3985), .C1(n183), .C2(n4019), .A(n1222), 
        .ZN(n1231) );
  OAI22_X1 U1163 ( .A1(n192), .A2(n1224), .B1(n189), .B2(n1223), .ZN(n1225) );
  AOI221_X1 U1164 ( .B1(n198), .B2(n4125), .C1(n195), .C2(n4160), .A(n1225), 
        .ZN(n1230) );
  OAI22_X1 U1165 ( .A1(n204), .A2(n1227), .B1(n201), .B2(n1226), .ZN(n1228) );
  AOI221_X1 U1166 ( .B1(n210), .B2(n4265), .C1(n207), .C2(n4305), .A(n1228), 
        .ZN(n1229) );
  NAND4_X1 U1167 ( .A1(n1232), .A2(n1231), .A3(n1230), .A4(n1229), .ZN(n1250)
         );
  OAI22_X1 U1168 ( .A1(n216), .A2(n1234), .B1(n213), .B2(n1233), .ZN(n1235) );
  AOI221_X1 U1169 ( .B1(n222), .B2(n2280), .C1(n219), .C2(n2314), .A(n1235), 
        .ZN(n1248) );
  OAI22_X1 U1170 ( .A1(n228), .A2(n1237), .B1(n225), .B2(n1236), .ZN(n1238) );
  AOI221_X1 U1171 ( .B1(n234), .B2(n2416), .C1(n231), .C2(n2454), .A(n1238), 
        .ZN(n1247) );
  OAI22_X1 U1172 ( .A1(n240), .A2(n1240), .B1(n237), .B2(n1239), .ZN(n1241) );
  AOI221_X1 U1173 ( .B1(n246), .B2(n2488), .C1(n243), .C2(n2522), .A(n1241), 
        .ZN(n1246) );
  OAI22_X1 U1174 ( .A1(n252), .A2(n1243), .B1(n249), .B2(n1242), .ZN(n1244) );
  AOI221_X1 U1175 ( .B1(n258), .B2(n3712), .C1(n255), .C2(n3746), .A(n1244), 
        .ZN(n1245) );
  NAND4_X1 U1176 ( .A1(n1248), .A2(n1247), .A3(n1246), .A4(n1245), .ZN(n1249)
         );
  OAI21_X1 U1177 ( .B1(n1250), .B2(n1249), .A(n261), .ZN(n1251) );
  OAI21_X1 U1178 ( .B1(n264), .B2(n1252), .A(n1251), .ZN(n2564) );
  OAI22_X1 U1179 ( .A1(n168), .A2(n1254), .B1(n165), .B2(n1253), .ZN(n1255) );
  AOI221_X1 U1180 ( .B1(n174), .B2(n3850), .C1(n171), .C2(n3884), .A(n1255), 
        .ZN(n1268) );
  OAI22_X1 U1181 ( .A1(n180), .A2(n1257), .B1(n177), .B2(n1256), .ZN(n1258) );
  AOI221_X1 U1182 ( .B1(n186), .B2(n3986), .C1(n183), .C2(n4020), .A(n1258), 
        .ZN(n1267) );
  OAI22_X1 U1183 ( .A1(n192), .A2(n1260), .B1(n189), .B2(n1259), .ZN(n1261) );
  AOI221_X1 U1184 ( .B1(n198), .B2(n4126), .C1(n195), .C2(n4161), .A(n1261), 
        .ZN(n1266) );
  OAI22_X1 U1185 ( .A1(n204), .A2(n1263), .B1(n201), .B2(n1262), .ZN(n1264) );
  AOI221_X1 U1186 ( .B1(n210), .B2(n4266), .C1(n207), .C2(n4307), .A(n1264), 
        .ZN(n1265) );
  NAND4_X1 U1187 ( .A1(n1268), .A2(n1267), .A3(n1266), .A4(n1265), .ZN(n1286)
         );
  OAI22_X1 U1188 ( .A1(n216), .A2(n1270), .B1(n213), .B2(n1269), .ZN(n1271) );
  AOI221_X1 U1189 ( .B1(n222), .B2(n2281), .C1(n219), .C2(n2315), .A(n1271), 
        .ZN(n1284) );
  OAI22_X1 U1190 ( .A1(n228), .A2(n1273), .B1(n225), .B2(n1272), .ZN(n1274) );
  AOI221_X1 U1191 ( .B1(n234), .B2(n2417), .C1(n231), .C2(n2455), .A(n1274), 
        .ZN(n1283) );
  OAI22_X1 U1192 ( .A1(n240), .A2(n1276), .B1(n237), .B2(n1275), .ZN(n1277) );
  AOI221_X1 U1193 ( .B1(n246), .B2(n2489), .C1(n243), .C2(n2523), .A(n1277), 
        .ZN(n1282) );
  OAI22_X1 U1194 ( .A1(n252), .A2(n1279), .B1(n249), .B2(n1278), .ZN(n1280) );
  AOI221_X1 U1195 ( .B1(n258), .B2(n3713), .C1(n255), .C2(n3747), .A(n1280), 
        .ZN(n1281) );
  NAND4_X1 U1196 ( .A1(n1284), .A2(n1283), .A3(n1282), .A4(n1281), .ZN(n1285)
         );
  OAI21_X1 U1197 ( .B1(n1286), .B2(n1285), .A(n261), .ZN(n1287) );
  OAI21_X1 U1198 ( .B1(n264), .B2(n1288), .A(n1287), .ZN(n2565) );
  OAI22_X1 U1199 ( .A1(n168), .A2(n1290), .B1(n165), .B2(n1289), .ZN(n1291) );
  AOI221_X1 U1200 ( .B1(n174), .B2(n3851), .C1(n171), .C2(n3885), .A(n1291), 
        .ZN(n1304) );
  OAI22_X1 U1201 ( .A1(n180), .A2(n1293), .B1(n177), .B2(n1292), .ZN(n1294) );
  AOI221_X1 U1202 ( .B1(n186), .B2(n3987), .C1(n183), .C2(n4021), .A(n1294), 
        .ZN(n1303) );
  OAI22_X1 U1203 ( .A1(n192), .A2(n1296), .B1(n189), .B2(n1295), .ZN(n1297) );
  AOI221_X1 U1204 ( .B1(n198), .B2(n4127), .C1(n195), .C2(n4162), .A(n1297), 
        .ZN(n1302) );
  OAI22_X1 U1205 ( .A1(n204), .A2(n1299), .B1(n201), .B2(n1298), .ZN(n1300) );
  AOI221_X1 U1206 ( .B1(n210), .B2(n4267), .C1(n207), .C2(n4309), .A(n1300), 
        .ZN(n1301) );
  NAND4_X1 U1207 ( .A1(n1304), .A2(n1303), .A3(n1302), .A4(n1301), .ZN(n1322)
         );
  OAI22_X1 U1208 ( .A1(n216), .A2(n1306), .B1(n213), .B2(n1305), .ZN(n1307) );
  AOI221_X1 U1209 ( .B1(n222), .B2(n2282), .C1(n219), .C2(n2316), .A(n1307), 
        .ZN(n1320) );
  OAI22_X1 U1210 ( .A1(n228), .A2(n1309), .B1(n225), .B2(n1308), .ZN(n1310) );
  AOI221_X1 U1211 ( .B1(n234), .B2(n2418), .C1(n231), .C2(n2456), .A(n1310), 
        .ZN(n1319) );
  OAI22_X1 U1212 ( .A1(n240), .A2(n1312), .B1(n237), .B2(n1311), .ZN(n1313) );
  AOI221_X1 U1213 ( .B1(n246), .B2(n2490), .C1(n243), .C2(n2524), .A(n1313), 
        .ZN(n1318) );
  OAI22_X1 U1214 ( .A1(n252), .A2(n1315), .B1(n249), .B2(n1314), .ZN(n1316) );
  AOI221_X1 U1215 ( .B1(n258), .B2(n3714), .C1(n255), .C2(n3748), .A(n1316), 
        .ZN(n1317) );
  NAND4_X1 U1216 ( .A1(n1320), .A2(n1319), .A3(n1318), .A4(n1317), .ZN(n1321)
         );
  OAI21_X1 U1217 ( .B1(n1322), .B2(n1321), .A(n261), .ZN(n1323) );
  OAI21_X1 U1218 ( .B1(n264), .B2(n1324), .A(n1323), .ZN(n2566) );
  OAI22_X1 U1219 ( .A1(n168), .A2(n1326), .B1(n165), .B2(n1325), .ZN(n1327) );
  AOI221_X1 U1220 ( .B1(n174), .B2(n3852), .C1(n171), .C2(n3886), .A(n1327), 
        .ZN(n1340) );
  OAI22_X1 U1221 ( .A1(n180), .A2(n1329), .B1(n177), .B2(n1328), .ZN(n1330) );
  AOI221_X1 U1222 ( .B1(n186), .B2(n3988), .C1(n183), .C2(n4022), .A(n1330), 
        .ZN(n1339) );
  OAI22_X1 U1223 ( .A1(n192), .A2(n1332), .B1(n189), .B2(n1331), .ZN(n1333) );
  AOI221_X1 U1224 ( .B1(n198), .B2(n4128), .C1(n195), .C2(n4163), .A(n1333), 
        .ZN(n1338) );
  OAI22_X1 U1225 ( .A1(n204), .A2(n1335), .B1(n201), .B2(n1334), .ZN(n1336) );
  AOI221_X1 U1226 ( .B1(n210), .B2(n4268), .C1(n207), .C2(n4311), .A(n1336), 
        .ZN(n1337) );
  NAND4_X1 U1227 ( .A1(n1340), .A2(n1339), .A3(n1338), .A4(n1337), .ZN(n1358)
         );
  OAI22_X1 U1228 ( .A1(n216), .A2(n1342), .B1(n213), .B2(n1341), .ZN(n1343) );
  AOI221_X1 U1229 ( .B1(n222), .B2(n2283), .C1(n219), .C2(n2317), .A(n1343), 
        .ZN(n1356) );
  OAI22_X1 U1230 ( .A1(n228), .A2(n1345), .B1(n225), .B2(n1344), .ZN(n1346) );
  AOI221_X1 U1231 ( .B1(n234), .B2(n2419), .C1(n231), .C2(n2457), .A(n1346), 
        .ZN(n1355) );
  OAI22_X1 U1232 ( .A1(n240), .A2(n1348), .B1(n237), .B2(n1347), .ZN(n1349) );
  AOI221_X1 U1233 ( .B1(n246), .B2(n2491), .C1(n243), .C2(n2525), .A(n1349), 
        .ZN(n1354) );
  OAI22_X1 U1234 ( .A1(n252), .A2(n1351), .B1(n249), .B2(n1350), .ZN(n1352) );
  AOI221_X1 U1235 ( .B1(n258), .B2(n3715), .C1(n255), .C2(n3749), .A(n1352), 
        .ZN(n1353) );
  NAND4_X1 U1236 ( .A1(n1356), .A2(n1355), .A3(n1354), .A4(n1353), .ZN(n1357)
         );
  OAI21_X1 U1237 ( .B1(n1358), .B2(n1357), .A(n261), .ZN(n1359) );
  OAI21_X1 U1238 ( .B1(n264), .B2(n1360), .A(n1359), .ZN(n2567) );
  OAI22_X1 U1239 ( .A1(n168), .A2(n1362), .B1(n165), .B2(n1361), .ZN(n1363) );
  AOI221_X1 U1240 ( .B1(n174), .B2(n3853), .C1(n171), .C2(n3887), .A(n1363), 
        .ZN(n1376) );
  OAI22_X1 U1241 ( .A1(n180), .A2(n1365), .B1(n177), .B2(n1364), .ZN(n1366) );
  AOI221_X1 U1242 ( .B1(n186), .B2(n3989), .C1(n183), .C2(n4023), .A(n1366), 
        .ZN(n1375) );
  OAI22_X1 U1243 ( .A1(n192), .A2(n1368), .B1(n189), .B2(n1367), .ZN(n1369) );
  AOI221_X1 U1244 ( .B1(n198), .B2(n4129), .C1(n195), .C2(n4164), .A(n1369), 
        .ZN(n1374) );
  OAI22_X1 U1245 ( .A1(n204), .A2(n1371), .B1(n201), .B2(n1370), .ZN(n1372) );
  AOI221_X1 U1246 ( .B1(n210), .B2(n4269), .C1(n207), .C2(n4313), .A(n1372), 
        .ZN(n1373) );
  NAND4_X1 U1247 ( .A1(n1376), .A2(n1375), .A3(n1374), .A4(n1373), .ZN(n1394)
         );
  OAI22_X1 U1248 ( .A1(n216), .A2(n1378), .B1(n213), .B2(n1377), .ZN(n1379) );
  AOI221_X1 U1249 ( .B1(n222), .B2(n2284), .C1(n219), .C2(n2318), .A(n1379), 
        .ZN(n1392) );
  OAI22_X1 U1250 ( .A1(n228), .A2(n1381), .B1(n225), .B2(n1380), .ZN(n1382) );
  AOI221_X1 U1251 ( .B1(n234), .B2(n2420), .C1(n231), .C2(n2458), .A(n1382), 
        .ZN(n1391) );
  OAI22_X1 U1252 ( .A1(n240), .A2(n1384), .B1(n237), .B2(n1383), .ZN(n1385) );
  AOI221_X1 U1253 ( .B1(n246), .B2(n2492), .C1(n243), .C2(n2526), .A(n1385), 
        .ZN(n1390) );
  OAI22_X1 U1254 ( .A1(n252), .A2(n1387), .B1(n249), .B2(n1386), .ZN(n1388) );
  AOI221_X1 U1255 ( .B1(n258), .B2(n3716), .C1(n255), .C2(n3750), .A(n1388), 
        .ZN(n1389) );
  NAND4_X1 U1256 ( .A1(n1392), .A2(n1391), .A3(n1390), .A4(n1389), .ZN(n1393)
         );
  OAI21_X1 U1257 ( .B1(n1394), .B2(n1393), .A(n261), .ZN(n1395) );
  OAI21_X1 U1258 ( .B1(n264), .B2(n1396), .A(n1395), .ZN(n2568) );
  OAI22_X1 U1259 ( .A1(n168), .A2(n1398), .B1(n165), .B2(n1397), .ZN(n1399) );
  AOI221_X1 U1260 ( .B1(n174), .B2(n3854), .C1(n171), .C2(n3888), .A(n1399), 
        .ZN(n1412) );
  OAI22_X1 U1261 ( .A1(n180), .A2(n1401), .B1(n177), .B2(n1400), .ZN(n1402) );
  AOI221_X1 U1262 ( .B1(n186), .B2(n3990), .C1(n183), .C2(n4024), .A(n1402), 
        .ZN(n1411) );
  OAI22_X1 U1263 ( .A1(n192), .A2(n1404), .B1(n189), .B2(n1403), .ZN(n1405) );
  AOI221_X1 U1264 ( .B1(n198), .B2(n4130), .C1(n195), .C2(n4165), .A(n1405), 
        .ZN(n1410) );
  OAI22_X1 U1265 ( .A1(n204), .A2(n1407), .B1(n201), .B2(n1406), .ZN(n1408) );
  AOI221_X1 U1266 ( .B1(n210), .B2(n4270), .C1(n207), .C2(n4315), .A(n1408), 
        .ZN(n1409) );
  NAND4_X1 U1267 ( .A1(n1412), .A2(n1411), .A3(n1410), .A4(n1409), .ZN(n1430)
         );
  OAI22_X1 U1268 ( .A1(n216), .A2(n1414), .B1(n213), .B2(n1413), .ZN(n1415) );
  AOI221_X1 U1269 ( .B1(n222), .B2(n2285), .C1(n219), .C2(n2319), .A(n1415), 
        .ZN(n1428) );
  OAI22_X1 U1270 ( .A1(n228), .A2(n1417), .B1(n225), .B2(n1416), .ZN(n1418) );
  AOI221_X1 U1271 ( .B1(n234), .B2(n2421), .C1(n231), .C2(n2459), .A(n1418), 
        .ZN(n1427) );
  OAI22_X1 U1272 ( .A1(n240), .A2(n1420), .B1(n237), .B2(n1419), .ZN(n1421) );
  AOI221_X1 U1273 ( .B1(n246), .B2(n2493), .C1(n243), .C2(n3615), .A(n1421), 
        .ZN(n1426) );
  OAI22_X1 U1274 ( .A1(n252), .A2(n1423), .B1(n249), .B2(n1422), .ZN(n1424) );
  AOI221_X1 U1275 ( .B1(n258), .B2(n3717), .C1(n255), .C2(n3751), .A(n1424), 
        .ZN(n1425) );
  NAND4_X1 U1276 ( .A1(n1428), .A2(n1427), .A3(n1426), .A4(n1425), .ZN(n1429)
         );
  OAI21_X1 U1277 ( .B1(n1430), .B2(n1429), .A(n261), .ZN(n1431) );
  OAI21_X1 U1278 ( .B1(n264), .B2(n1432), .A(n1431), .ZN(n2569) );
  OAI22_X1 U1279 ( .A1(n168), .A2(n1434), .B1(n165), .B2(n1433), .ZN(n1435) );
  AOI221_X1 U1280 ( .B1(n174), .B2(n3855), .C1(n171), .C2(n3889), .A(n1435), 
        .ZN(n1448) );
  OAI22_X1 U1281 ( .A1(n180), .A2(n1437), .B1(n177), .B2(n1436), .ZN(n1438) );
  AOI221_X1 U1282 ( .B1(n186), .B2(n3991), .C1(n183), .C2(n4025), .A(n1438), 
        .ZN(n1447) );
  OAI22_X1 U1283 ( .A1(n192), .A2(n1440), .B1(n189), .B2(n1439), .ZN(n1441) );
  AOI221_X1 U1284 ( .B1(n198), .B2(n4131), .C1(n195), .C2(n4166), .A(n1441), 
        .ZN(n1446) );
  OAI22_X1 U1285 ( .A1(n204), .A2(n1443), .B1(n201), .B2(n1442), .ZN(n1444) );
  AOI221_X1 U1286 ( .B1(n210), .B2(n4271), .C1(n207), .C2(n4317), .A(n1444), 
        .ZN(n1445) );
  NAND4_X1 U1287 ( .A1(n1448), .A2(n1447), .A3(n1446), .A4(n1445), .ZN(n1466)
         );
  OAI22_X1 U1288 ( .A1(n216), .A2(n1450), .B1(n213), .B2(n1449), .ZN(n1451) );
  AOI221_X1 U1289 ( .B1(n222), .B2(n2286), .C1(n219), .C2(n2320), .A(n1451), 
        .ZN(n1464) );
  OAI22_X1 U1290 ( .A1(n228), .A2(n1453), .B1(n225), .B2(n1452), .ZN(n1454) );
  AOI221_X1 U1291 ( .B1(n234), .B2(n2422), .C1(n231), .C2(n2460), .A(n1454), 
        .ZN(n1463) );
  OAI22_X1 U1292 ( .A1(n240), .A2(n1456), .B1(n237), .B2(n1455), .ZN(n1457) );
  AOI221_X1 U1293 ( .B1(n246), .B2(n2494), .C1(n243), .C2(n3616), .A(n1457), 
        .ZN(n1462) );
  OAI22_X1 U1294 ( .A1(n252), .A2(n1459), .B1(n249), .B2(n1458), .ZN(n1460) );
  AOI221_X1 U1295 ( .B1(n258), .B2(n3718), .C1(n255), .C2(n3752), .A(n1460), 
        .ZN(n1461) );
  NAND4_X1 U1296 ( .A1(n1464), .A2(n1463), .A3(n1462), .A4(n1461), .ZN(n1465)
         );
  OAI21_X1 U1297 ( .B1(n1466), .B2(n1465), .A(n261), .ZN(n1467) );
  OAI21_X1 U1298 ( .B1(n265), .B2(n1468), .A(n1467), .ZN(n2570) );
  OAI22_X1 U1299 ( .A1(n169), .A2(n1470), .B1(n166), .B2(n1469), .ZN(n1471) );
  AOI221_X1 U1300 ( .B1(n175), .B2(n3856), .C1(n172), .C2(n3890), .A(n1471), 
        .ZN(n1484) );
  OAI22_X1 U1301 ( .A1(n181), .A2(n1473), .B1(n178), .B2(n1472), .ZN(n1474) );
  AOI221_X1 U1302 ( .B1(n187), .B2(n3992), .C1(n184), .C2(n4026), .A(n1474), 
        .ZN(n1483) );
  OAI22_X1 U1303 ( .A1(n193), .A2(n1476), .B1(n190), .B2(n1475), .ZN(n1477) );
  AOI221_X1 U1304 ( .B1(n199), .B2(n4132), .C1(n196), .C2(n4167), .A(n1477), 
        .ZN(n1482) );
  OAI22_X1 U1305 ( .A1(n205), .A2(n1479), .B1(n202), .B2(n1478), .ZN(n1480) );
  AOI221_X1 U1306 ( .B1(n211), .B2(n4272), .C1(n208), .C2(n4319), .A(n1480), 
        .ZN(n1481) );
  NAND4_X1 U1307 ( .A1(n1484), .A2(n1483), .A3(n1482), .A4(n1481), .ZN(n1502)
         );
  OAI22_X1 U1308 ( .A1(n217), .A2(n1486), .B1(n214), .B2(n1485), .ZN(n1487) );
  AOI221_X1 U1309 ( .B1(n223), .B2(n2287), .C1(n220), .C2(n2321), .A(n1487), 
        .ZN(n1500) );
  OAI22_X1 U1310 ( .A1(n229), .A2(n1489), .B1(n226), .B2(n1488), .ZN(n1490) );
  AOI221_X1 U1311 ( .B1(n235), .B2(n2423), .C1(n232), .C2(n2461), .A(n1490), 
        .ZN(n1499) );
  OAI22_X1 U1312 ( .A1(n241), .A2(n1492), .B1(n238), .B2(n1491), .ZN(n1493) );
  AOI221_X1 U1313 ( .B1(n247), .B2(n2495), .C1(n244), .C2(n3617), .A(n1493), 
        .ZN(n1498) );
  OAI22_X1 U1314 ( .A1(n253), .A2(n1495), .B1(n250), .B2(n1494), .ZN(n1496) );
  AOI221_X1 U1315 ( .B1(n259), .B2(n3719), .C1(n256), .C2(n3753), .A(n1496), 
        .ZN(n1497) );
  NAND4_X1 U1316 ( .A1(n1500), .A2(n1499), .A3(n1498), .A4(n1497), .ZN(n1501)
         );
  OAI21_X1 U1317 ( .B1(n1502), .B2(n1501), .A(n262), .ZN(n1503) );
  OAI21_X1 U1318 ( .B1(n265), .B2(n1504), .A(n1503), .ZN(n2571) );
  OAI22_X1 U1319 ( .A1(n169), .A2(n1506), .B1(n166), .B2(n1505), .ZN(n1507) );
  AOI221_X1 U1320 ( .B1(n175), .B2(n3857), .C1(n172), .C2(n3891), .A(n1507), 
        .ZN(n1520) );
  OAI22_X1 U1321 ( .A1(n181), .A2(n1509), .B1(n178), .B2(n1508), .ZN(n1510) );
  AOI221_X1 U1322 ( .B1(n187), .B2(n3993), .C1(n184), .C2(n4027), .A(n1510), 
        .ZN(n1519) );
  OAI22_X1 U1323 ( .A1(n193), .A2(n1512), .B1(n190), .B2(n1511), .ZN(n1513) );
  AOI221_X1 U1324 ( .B1(n199), .B2(n4133), .C1(n196), .C2(n4168), .A(n1513), 
        .ZN(n1518) );
  OAI22_X1 U1325 ( .A1(n205), .A2(n1515), .B1(n202), .B2(n1514), .ZN(n1516) );
  AOI221_X1 U1326 ( .B1(n211), .B2(n4273), .C1(n208), .C2(n4321), .A(n1516), 
        .ZN(n1517) );
  NAND4_X1 U1327 ( .A1(n1520), .A2(n1519), .A3(n1518), .A4(n1517), .ZN(n1538)
         );
  OAI22_X1 U1328 ( .A1(n217), .A2(n1522), .B1(n214), .B2(n1521), .ZN(n1523) );
  AOI221_X1 U1329 ( .B1(n223), .B2(n2288), .C1(n220), .C2(n2322), .A(n1523), 
        .ZN(n1536) );
  OAI22_X1 U1330 ( .A1(n229), .A2(n1525), .B1(n226), .B2(n1524), .ZN(n1526) );
  AOI221_X1 U1331 ( .B1(n235), .B2(n2424), .C1(n232), .C2(n2462), .A(n1526), 
        .ZN(n1535) );
  OAI22_X1 U1332 ( .A1(n241), .A2(n1528), .B1(n238), .B2(n1527), .ZN(n1529) );
  AOI221_X1 U1333 ( .B1(n247), .B2(n2496), .C1(n244), .C2(n3618), .A(n1529), 
        .ZN(n1534) );
  OAI22_X1 U1334 ( .A1(n253), .A2(n1531), .B1(n250), .B2(n1530), .ZN(n1532) );
  AOI221_X1 U1335 ( .B1(n259), .B2(n3720), .C1(n256), .C2(n3754), .A(n1532), 
        .ZN(n1533) );
  NAND4_X1 U1336 ( .A1(n1536), .A2(n1535), .A3(n1534), .A4(n1533), .ZN(n1537)
         );
  OAI21_X1 U1337 ( .B1(n1538), .B2(n1537), .A(n262), .ZN(n1539) );
  OAI21_X1 U1338 ( .B1(n265), .B2(n1540), .A(n1539), .ZN(n2572) );
  OAI22_X1 U1339 ( .A1(n169), .A2(n1542), .B1(n166), .B2(n1541), .ZN(n1543) );
  AOI221_X1 U1340 ( .B1(n175), .B2(n3858), .C1(n172), .C2(n3892), .A(n1543), 
        .ZN(n1556) );
  OAI22_X1 U1341 ( .A1(n181), .A2(n1545), .B1(n178), .B2(n1544), .ZN(n1546) );
  AOI221_X1 U1342 ( .B1(n187), .B2(n3994), .C1(n184), .C2(n4028), .A(n1546), 
        .ZN(n1555) );
  OAI22_X1 U1343 ( .A1(n193), .A2(n1548), .B1(n190), .B2(n1547), .ZN(n1549) );
  AOI221_X1 U1344 ( .B1(n199), .B2(n4134), .C1(n196), .C2(n4169), .A(n1549), 
        .ZN(n1554) );
  OAI22_X1 U1345 ( .A1(n205), .A2(n1551), .B1(n202), .B2(n1550), .ZN(n1552) );
  AOI221_X1 U1346 ( .B1(n211), .B2(n4274), .C1(n208), .C2(n4323), .A(n1552), 
        .ZN(n1553) );
  NAND4_X1 U1347 ( .A1(n1556), .A2(n1555), .A3(n1554), .A4(n1553), .ZN(n1574)
         );
  OAI22_X1 U1348 ( .A1(n217), .A2(n1558), .B1(n214), .B2(n1557), .ZN(n1559) );
  AOI221_X1 U1349 ( .B1(n223), .B2(n2289), .C1(n220), .C2(n2323), .A(n1559), 
        .ZN(n1572) );
  OAI22_X1 U1350 ( .A1(n229), .A2(n1561), .B1(n226), .B2(n1560), .ZN(n1562) );
  AOI221_X1 U1351 ( .B1(n235), .B2(n2425), .C1(n232), .C2(n2463), .A(n1562), 
        .ZN(n1571) );
  OAI22_X1 U1352 ( .A1(n241), .A2(n1564), .B1(n238), .B2(n1563), .ZN(n1565) );
  AOI221_X1 U1353 ( .B1(n247), .B2(n2497), .C1(n244), .C2(n3619), .A(n1565), 
        .ZN(n1570) );
  OAI22_X1 U1354 ( .A1(n253), .A2(n1567), .B1(n250), .B2(n1566), .ZN(n1568) );
  AOI221_X1 U1355 ( .B1(n259), .B2(n3721), .C1(n256), .C2(n3755), .A(n1568), 
        .ZN(n1569) );
  NAND4_X1 U1356 ( .A1(n1572), .A2(n1571), .A3(n1570), .A4(n1569), .ZN(n1573)
         );
  OAI21_X1 U1357 ( .B1(n1574), .B2(n1573), .A(n262), .ZN(n1575) );
  OAI21_X1 U1358 ( .B1(n265), .B2(n1576), .A(n1575), .ZN(n2573) );
  OAI22_X1 U1359 ( .A1(n169), .A2(n1578), .B1(n166), .B2(n1577), .ZN(n1579) );
  AOI221_X1 U1360 ( .B1(n175), .B2(n3859), .C1(n172), .C2(n3893), .A(n1579), 
        .ZN(n1592) );
  OAI22_X1 U1361 ( .A1(n181), .A2(n1581), .B1(n178), .B2(n1580), .ZN(n1582) );
  AOI221_X1 U1362 ( .B1(n187), .B2(n3995), .C1(n184), .C2(n4029), .A(n1582), 
        .ZN(n1591) );
  OAI22_X1 U1363 ( .A1(n193), .A2(n1584), .B1(n190), .B2(n1583), .ZN(n1585) );
  AOI221_X1 U1364 ( .B1(n199), .B2(n4135), .C1(n196), .C2(n4170), .A(n1585), 
        .ZN(n1590) );
  OAI22_X1 U1365 ( .A1(n205), .A2(n1587), .B1(n202), .B2(n1586), .ZN(n1588) );
  AOI221_X1 U1366 ( .B1(n211), .B2(n4275), .C1(n208), .C2(n4325), .A(n1588), 
        .ZN(n1589) );
  NAND4_X1 U1367 ( .A1(n1592), .A2(n1591), .A3(n1590), .A4(n1589), .ZN(n1610)
         );
  OAI22_X1 U1368 ( .A1(n217), .A2(n1594), .B1(n214), .B2(n1593), .ZN(n1595) );
  AOI221_X1 U1369 ( .B1(n223), .B2(n2290), .C1(n220), .C2(n2324), .A(n1595), 
        .ZN(n1608) );
  OAI22_X1 U1370 ( .A1(n229), .A2(n1597), .B1(n226), .B2(n1596), .ZN(n1598) );
  AOI221_X1 U1371 ( .B1(n235), .B2(n2426), .C1(n232), .C2(n2464), .A(n1598), 
        .ZN(n1607) );
  OAI22_X1 U1372 ( .A1(n241), .A2(n1600), .B1(n238), .B2(n1599), .ZN(n1601) );
  AOI221_X1 U1373 ( .B1(n247), .B2(n2498), .C1(n244), .C2(n3620), .A(n1601), 
        .ZN(n1606) );
  OAI22_X1 U1374 ( .A1(n253), .A2(n1603), .B1(n250), .B2(n1602), .ZN(n1604) );
  AOI221_X1 U1375 ( .B1(n259), .B2(n3722), .C1(n256), .C2(n3756), .A(n1604), 
        .ZN(n1605) );
  NAND4_X1 U1376 ( .A1(n1608), .A2(n1607), .A3(n1606), .A4(n1605), .ZN(n1609)
         );
  OAI21_X1 U1377 ( .B1(n1610), .B2(n1609), .A(n262), .ZN(n1611) );
  OAI21_X1 U1378 ( .B1(n265), .B2(n1612), .A(n1611), .ZN(n2574) );
  OAI22_X1 U1379 ( .A1(n169), .A2(n1614), .B1(n166), .B2(n1613), .ZN(n1615) );
  AOI221_X1 U1380 ( .B1(n175), .B2(n3860), .C1(n172), .C2(n3894), .A(n1615), 
        .ZN(n1628) );
  OAI22_X1 U1381 ( .A1(n181), .A2(n1617), .B1(n178), .B2(n1616), .ZN(n1618) );
  AOI221_X1 U1382 ( .B1(n187), .B2(n3996), .C1(n184), .C2(n4030), .A(n1618), 
        .ZN(n1627) );
  OAI22_X1 U1383 ( .A1(n193), .A2(n1620), .B1(n190), .B2(n1619), .ZN(n1621) );
  AOI221_X1 U1384 ( .B1(n199), .B2(n4136), .C1(n196), .C2(n4171), .A(n1621), 
        .ZN(n1626) );
  OAI22_X1 U1385 ( .A1(n205), .A2(n1623), .B1(n202), .B2(n1622), .ZN(n1624) );
  AOI221_X1 U1386 ( .B1(n211), .B2(n4276), .C1(n208), .C2(n4327), .A(n1624), 
        .ZN(n1625) );
  NAND4_X1 U1387 ( .A1(n1628), .A2(n1627), .A3(n1626), .A4(n1625), .ZN(n1646)
         );
  OAI22_X1 U1388 ( .A1(n217), .A2(n1630), .B1(n214), .B2(n1629), .ZN(n1631) );
  AOI221_X1 U1389 ( .B1(n223), .B2(n2291), .C1(n220), .C2(n2325), .A(n1631), 
        .ZN(n1644) );
  OAI22_X1 U1390 ( .A1(n229), .A2(n1633), .B1(n226), .B2(n1632), .ZN(n1634) );
  AOI221_X1 U1391 ( .B1(n235), .B2(n2427), .C1(n232), .C2(n2465), .A(n1634), 
        .ZN(n1643) );
  OAI22_X1 U1392 ( .A1(n241), .A2(n1636), .B1(n238), .B2(n1635), .ZN(n1637) );
  AOI221_X1 U1393 ( .B1(n247), .B2(n2499), .C1(n244), .C2(n3621), .A(n1637), 
        .ZN(n1642) );
  OAI22_X1 U1394 ( .A1(n253), .A2(n1639), .B1(n250), .B2(n1638), .ZN(n1640) );
  AOI221_X1 U1395 ( .B1(n259), .B2(n3723), .C1(n256), .C2(n3757), .A(n1640), 
        .ZN(n1641) );
  NAND4_X1 U1396 ( .A1(n1644), .A2(n1643), .A3(n1642), .A4(n1641), .ZN(n1645)
         );
  OAI21_X1 U1397 ( .B1(n1646), .B2(n1645), .A(n262), .ZN(n1647) );
  OAI21_X1 U1398 ( .B1(n265), .B2(n1648), .A(n1647), .ZN(n2575) );
  OAI22_X1 U1399 ( .A1(n169), .A2(n1650), .B1(n166), .B2(n1649), .ZN(n1651) );
  AOI221_X1 U1400 ( .B1(n175), .B2(n3861), .C1(n172), .C2(n3895), .A(n1651), 
        .ZN(n1664) );
  OAI22_X1 U1401 ( .A1(n181), .A2(n1653), .B1(n178), .B2(n1652), .ZN(n1654) );
  AOI221_X1 U1402 ( .B1(n187), .B2(n3997), .C1(n184), .C2(n4031), .A(n1654), 
        .ZN(n1663) );
  OAI22_X1 U1403 ( .A1(n193), .A2(n1656), .B1(n190), .B2(n1655), .ZN(n1657) );
  AOI221_X1 U1404 ( .B1(n199), .B2(n4137), .C1(n196), .C2(n4172), .A(n1657), 
        .ZN(n1662) );
  OAI22_X1 U1405 ( .A1(n205), .A2(n1659), .B1(n202), .B2(n1658), .ZN(n1660) );
  AOI221_X1 U1406 ( .B1(n211), .B2(n4277), .C1(n208), .C2(n4329), .A(n1660), 
        .ZN(n1661) );
  NAND4_X1 U1407 ( .A1(n1664), .A2(n1663), .A3(n1662), .A4(n1661), .ZN(n1682)
         );
  OAI22_X1 U1408 ( .A1(n217), .A2(n1666), .B1(n214), .B2(n1665), .ZN(n1667) );
  AOI221_X1 U1409 ( .B1(n223), .B2(n2292), .C1(n220), .C2(n2326), .A(n1667), 
        .ZN(n1680) );
  OAI22_X1 U1410 ( .A1(n229), .A2(n1669), .B1(n226), .B2(n1668), .ZN(n1670) );
  AOI221_X1 U1411 ( .B1(n235), .B2(n2428), .C1(n232), .C2(n2466), .A(n1670), 
        .ZN(n1679) );
  OAI22_X1 U1412 ( .A1(n241), .A2(n1672), .B1(n238), .B2(n1671), .ZN(n1673) );
  AOI221_X1 U1413 ( .B1(n247), .B2(n2500), .C1(n244), .C2(n3622), .A(n1673), 
        .ZN(n1678) );
  OAI22_X1 U1414 ( .A1(n253), .A2(n1675), .B1(n250), .B2(n1674), .ZN(n1676) );
  AOI221_X1 U1415 ( .B1(n259), .B2(n3724), .C1(n256), .C2(n3758), .A(n1676), 
        .ZN(n1677) );
  NAND4_X1 U1416 ( .A1(n1680), .A2(n1679), .A3(n1678), .A4(n1677), .ZN(n1681)
         );
  OAI21_X1 U1417 ( .B1(n1682), .B2(n1681), .A(n262), .ZN(n1683) );
  OAI21_X1 U1418 ( .B1(n265), .B2(n1684), .A(n1683), .ZN(n2576) );
  OAI22_X1 U1419 ( .A1(n169), .A2(n1686), .B1(n166), .B2(n1685), .ZN(n1687) );
  AOI221_X1 U1420 ( .B1(n175), .B2(n3862), .C1(n172), .C2(n3896), .A(n1687), 
        .ZN(n1700) );
  OAI22_X1 U1421 ( .A1(n181), .A2(n1689), .B1(n178), .B2(n1688), .ZN(n1690) );
  AOI221_X1 U1422 ( .B1(n187), .B2(n3998), .C1(n184), .C2(n4032), .A(n1690), 
        .ZN(n1699) );
  OAI22_X1 U1423 ( .A1(n193), .A2(n1692), .B1(n190), .B2(n1691), .ZN(n1693) );
  AOI221_X1 U1424 ( .B1(n199), .B2(n4138), .C1(n196), .C2(n4173), .A(n1693), 
        .ZN(n1698) );
  OAI22_X1 U1425 ( .A1(n205), .A2(n1695), .B1(n202), .B2(n1694), .ZN(n1696) );
  AOI221_X1 U1426 ( .B1(n211), .B2(n4278), .C1(n208), .C2(n4331), .A(n1696), 
        .ZN(n1697) );
  NAND4_X1 U1427 ( .A1(n1700), .A2(n1699), .A3(n1698), .A4(n1697), .ZN(n1718)
         );
  OAI22_X1 U1428 ( .A1(n217), .A2(n1702), .B1(n214), .B2(n1701), .ZN(n1703) );
  AOI221_X1 U1429 ( .B1(n223), .B2(n2293), .C1(n220), .C2(n2327), .A(n1703), 
        .ZN(n1716) );
  OAI22_X1 U1430 ( .A1(n229), .A2(n1705), .B1(n226), .B2(n1704), .ZN(n1706) );
  AOI221_X1 U1431 ( .B1(n235), .B2(n2429), .C1(n232), .C2(n2467), .A(n1706), 
        .ZN(n1715) );
  OAI22_X1 U1432 ( .A1(n241), .A2(n1708), .B1(n238), .B2(n1707), .ZN(n1709) );
  AOI221_X1 U1433 ( .B1(n247), .B2(n2501), .C1(n244), .C2(n3623), .A(n1709), 
        .ZN(n1714) );
  OAI22_X1 U1434 ( .A1(n253), .A2(n1711), .B1(n250), .B2(n1710), .ZN(n1712) );
  AOI221_X1 U1435 ( .B1(n259), .B2(n3725), .C1(n256), .C2(n3759), .A(n1712), 
        .ZN(n1713) );
  NAND4_X1 U1436 ( .A1(n1716), .A2(n1715), .A3(n1714), .A4(n1713), .ZN(n1717)
         );
  OAI21_X1 U1437 ( .B1(n1718), .B2(n1717), .A(n262), .ZN(n1719) );
  OAI21_X1 U1438 ( .B1(n265), .B2(n1720), .A(n1719), .ZN(n2577) );
  OAI22_X1 U1439 ( .A1(n169), .A2(n1722), .B1(n166), .B2(n1721), .ZN(n1723) );
  AOI221_X1 U1440 ( .B1(n175), .B2(n3863), .C1(n172), .C2(n3897), .A(n1723), 
        .ZN(n1736) );
  OAI22_X1 U1441 ( .A1(n181), .A2(n1725), .B1(n178), .B2(n1724), .ZN(n1726) );
  AOI221_X1 U1442 ( .B1(n187), .B2(n3999), .C1(n184), .C2(n4033), .A(n1726), 
        .ZN(n1735) );
  OAI22_X1 U1443 ( .A1(n193), .A2(n1728), .B1(n190), .B2(n1727), .ZN(n1729) );
  AOI221_X1 U1444 ( .B1(n199), .B2(n4139), .C1(n196), .C2(n4174), .A(n1729), 
        .ZN(n1734) );
  OAI22_X1 U1445 ( .A1(n205), .A2(n1731), .B1(n202), .B2(n1730), .ZN(n1732) );
  AOI221_X1 U1446 ( .B1(n211), .B2(n4279), .C1(n208), .C2(n4333), .A(n1732), 
        .ZN(n1733) );
  NAND4_X1 U1447 ( .A1(n1736), .A2(n1735), .A3(n1734), .A4(n1733), .ZN(n1754)
         );
  OAI22_X1 U1448 ( .A1(n217), .A2(n1738), .B1(n214), .B2(n1737), .ZN(n1739) );
  AOI221_X1 U1449 ( .B1(n223), .B2(n2294), .C1(n220), .C2(n2328), .A(n1739), 
        .ZN(n1752) );
  OAI22_X1 U1450 ( .A1(n229), .A2(n1741), .B1(n226), .B2(n1740), .ZN(n1742) );
  AOI221_X1 U1451 ( .B1(n235), .B2(n2430), .C1(n232), .C2(n2468), .A(n1742), 
        .ZN(n1751) );
  OAI22_X1 U1452 ( .A1(n241), .A2(n1744), .B1(n238), .B2(n1743), .ZN(n1745) );
  AOI221_X1 U1453 ( .B1(n247), .B2(n2502), .C1(n244), .C2(n3624), .A(n1745), 
        .ZN(n1750) );
  OAI22_X1 U1454 ( .A1(n253), .A2(n1747), .B1(n250), .B2(n1746), .ZN(n1748) );
  AOI221_X1 U1455 ( .B1(n259), .B2(n3726), .C1(n256), .C2(n3760), .A(n1748), 
        .ZN(n1749) );
  NAND4_X1 U1456 ( .A1(n1752), .A2(n1751), .A3(n1750), .A4(n1749), .ZN(n1753)
         );
  OAI21_X1 U1457 ( .B1(n1754), .B2(n1753), .A(n262), .ZN(n1755) );
  OAI21_X1 U1458 ( .B1(n265), .B2(n1756), .A(n1755), .ZN(n2578) );
  OAI22_X1 U1459 ( .A1(n169), .A2(n1758), .B1(n166), .B2(n1757), .ZN(n1759) );
  AOI221_X1 U1460 ( .B1(n175), .B2(n3864), .C1(n172), .C2(n3898), .A(n1759), 
        .ZN(n1772) );
  OAI22_X1 U1461 ( .A1(n181), .A2(n1761), .B1(n178), .B2(n1760), .ZN(n1762) );
  AOI221_X1 U1462 ( .B1(n187), .B2(n4000), .C1(n184), .C2(n4034), .A(n1762), 
        .ZN(n1771) );
  OAI22_X1 U1463 ( .A1(n193), .A2(n1764), .B1(n190), .B2(n1763), .ZN(n1765) );
  AOI221_X1 U1464 ( .B1(n199), .B2(n4140), .C1(n196), .C2(n4175), .A(n1765), 
        .ZN(n1770) );
  OAI22_X1 U1465 ( .A1(n205), .A2(n1767), .B1(n202), .B2(n1766), .ZN(n1768) );
  AOI221_X1 U1466 ( .B1(n211), .B2(n4280), .C1(n208), .C2(n4335), .A(n1768), 
        .ZN(n1769) );
  NAND4_X1 U1467 ( .A1(n1772), .A2(n1771), .A3(n1770), .A4(n1769), .ZN(n1790)
         );
  OAI22_X1 U1468 ( .A1(n217), .A2(n1774), .B1(n214), .B2(n1773), .ZN(n1775) );
  AOI221_X1 U1469 ( .B1(n223), .B2(n2295), .C1(n220), .C2(n2329), .A(n1775), 
        .ZN(n1788) );
  OAI22_X1 U1470 ( .A1(n229), .A2(n1777), .B1(n226), .B2(n1776), .ZN(n1778) );
  AOI221_X1 U1471 ( .B1(n235), .B2(n2431), .C1(n232), .C2(n2469), .A(n1778), 
        .ZN(n1787) );
  OAI22_X1 U1472 ( .A1(n241), .A2(n1780), .B1(n238), .B2(n1779), .ZN(n1781) );
  AOI221_X1 U1473 ( .B1(n247), .B2(n2503), .C1(n244), .C2(n3625), .A(n1781), 
        .ZN(n1786) );
  OAI22_X1 U1474 ( .A1(n253), .A2(n1783), .B1(n250), .B2(n1782), .ZN(n1784) );
  AOI221_X1 U1475 ( .B1(n259), .B2(n3727), .C1(n256), .C2(n3761), .A(n1784), 
        .ZN(n1785) );
  NAND4_X1 U1476 ( .A1(n1788), .A2(n1787), .A3(n1786), .A4(n1785), .ZN(n1789)
         );
  OAI21_X1 U1477 ( .B1(n1790), .B2(n1789), .A(n262), .ZN(n1791) );
  OAI21_X1 U1478 ( .B1(n265), .B2(n1792), .A(n1791), .ZN(n2579) );
  OAI22_X1 U1479 ( .A1(n169), .A2(n1794), .B1(n166), .B2(n1793), .ZN(n1795) );
  AOI221_X1 U1480 ( .B1(n175), .B2(n3865), .C1(n172), .C2(n3899), .A(n1795), 
        .ZN(n1808) );
  OAI22_X1 U1481 ( .A1(n181), .A2(n1797), .B1(n178), .B2(n1796), .ZN(n1798) );
  AOI221_X1 U1482 ( .B1(n187), .B2(n4001), .C1(n184), .C2(n4035), .A(n1798), 
        .ZN(n1807) );
  OAI22_X1 U1483 ( .A1(n193), .A2(n1800), .B1(n190), .B2(n1799), .ZN(n1801) );
  AOI221_X1 U1484 ( .B1(n199), .B2(n4141), .C1(n196), .C2(n4176), .A(n1801), 
        .ZN(n1806) );
  OAI22_X1 U1485 ( .A1(n205), .A2(n1803), .B1(n202), .B2(n1802), .ZN(n1804) );
  AOI221_X1 U1486 ( .B1(n211), .B2(n4281), .C1(n208), .C2(n4337), .A(n1804), 
        .ZN(n1805) );
  NAND4_X1 U1487 ( .A1(n1808), .A2(n1807), .A3(n1806), .A4(n1805), .ZN(n1826)
         );
  OAI22_X1 U1488 ( .A1(n217), .A2(n1810), .B1(n214), .B2(n1809), .ZN(n1811) );
  AOI221_X1 U1489 ( .B1(n223), .B2(n2296), .C1(n220), .C2(n2330), .A(n1811), 
        .ZN(n1824) );
  OAI22_X1 U1490 ( .A1(n229), .A2(n1813), .B1(n226), .B2(n1812), .ZN(n1814) );
  AOI221_X1 U1491 ( .B1(n235), .B2(n2432), .C1(n232), .C2(n2470), .A(n1814), 
        .ZN(n1823) );
  OAI22_X1 U1492 ( .A1(n241), .A2(n1816), .B1(n238), .B2(n1815), .ZN(n1817) );
  AOI221_X1 U1493 ( .B1(n247), .B2(n2504), .C1(n244), .C2(n3626), .A(n1817), 
        .ZN(n1822) );
  OAI22_X1 U1494 ( .A1(n253), .A2(n1819), .B1(n250), .B2(n1818), .ZN(n1820) );
  AOI221_X1 U1495 ( .B1(n259), .B2(n3728), .C1(n256), .C2(n3762), .A(n1820), 
        .ZN(n1821) );
  NAND4_X1 U1496 ( .A1(n1824), .A2(n1823), .A3(n1822), .A4(n1821), .ZN(n1825)
         );
  OAI21_X1 U1497 ( .B1(n1826), .B2(n1825), .A(n262), .ZN(n1827) );
  OAI21_X1 U1498 ( .B1(n265), .B2(n1828), .A(n1827), .ZN(n2580) );
  OAI22_X1 U1499 ( .A1(n169), .A2(n1830), .B1(n166), .B2(n1829), .ZN(n1831) );
  AOI221_X1 U1500 ( .B1(n175), .B2(n3866), .C1(n172), .C2(n3900), .A(n1831), 
        .ZN(n1844) );
  OAI22_X1 U1501 ( .A1(n181), .A2(n1833), .B1(n178), .B2(n1832), .ZN(n1834) );
  AOI221_X1 U1502 ( .B1(n187), .B2(n4002), .C1(n184), .C2(n4036), .A(n1834), 
        .ZN(n1843) );
  OAI22_X1 U1503 ( .A1(n193), .A2(n1836), .B1(n190), .B2(n1835), .ZN(n1837) );
  AOI221_X1 U1504 ( .B1(n199), .B2(n4142), .C1(n196), .C2(n4177), .A(n1837), 
        .ZN(n1842) );
  OAI22_X1 U1505 ( .A1(n205), .A2(n1839), .B1(n202), .B2(n1838), .ZN(n1840) );
  AOI221_X1 U1506 ( .B1(n211), .B2(n4282), .C1(n208), .C2(n4339), .A(n1840), 
        .ZN(n1841) );
  NAND4_X1 U1507 ( .A1(n1844), .A2(n1843), .A3(n1842), .A4(n1841), .ZN(n1862)
         );
  OAI22_X1 U1508 ( .A1(n217), .A2(n1846), .B1(n214), .B2(n1845), .ZN(n1847) );
  AOI221_X1 U1509 ( .B1(n223), .B2(n2297), .C1(n220), .C2(n2331), .A(n1847), 
        .ZN(n1860) );
  OAI22_X1 U1510 ( .A1(n229), .A2(n1849), .B1(n226), .B2(n1848), .ZN(n1850) );
  AOI221_X1 U1511 ( .B1(n235), .B2(n2433), .C1(n232), .C2(n2471), .A(n1850), 
        .ZN(n1859) );
  OAI22_X1 U1512 ( .A1(n241), .A2(n1852), .B1(n238), .B2(n1851), .ZN(n1853) );
  AOI221_X1 U1513 ( .B1(n247), .B2(n2505), .C1(n244), .C2(n3627), .A(n1853), 
        .ZN(n1858) );
  OAI22_X1 U1514 ( .A1(n253), .A2(n1855), .B1(n250), .B2(n1854), .ZN(n1856) );
  AOI221_X1 U1515 ( .B1(n259), .B2(n3729), .C1(n256), .C2(n3763), .A(n1856), 
        .ZN(n1857) );
  NAND4_X1 U1516 ( .A1(n1860), .A2(n1859), .A3(n1858), .A4(n1857), .ZN(n1861)
         );
  OAI21_X1 U1517 ( .B1(n1862), .B2(n1861), .A(n262), .ZN(n1863) );
  OAI21_X1 U1518 ( .B1(n265), .B2(n1864), .A(n1863), .ZN(n2581) );
  OAI22_X1 U1519 ( .A1(n169), .A2(n1866), .B1(n166), .B2(n1865), .ZN(n1867) );
  AOI221_X1 U1520 ( .B1(n175), .B2(n3867), .C1(n172), .C2(n3901), .A(n1867), 
        .ZN(n1880) );
  OAI22_X1 U1521 ( .A1(n181), .A2(n1869), .B1(n178), .B2(n1868), .ZN(n1870) );
  AOI221_X1 U1522 ( .B1(n187), .B2(n4003), .C1(n184), .C2(n4037), .A(n1870), 
        .ZN(n1879) );
  OAI22_X1 U1523 ( .A1(n193), .A2(n1872), .B1(n190), .B2(n1871), .ZN(n1873) );
  AOI221_X1 U1524 ( .B1(n199), .B2(n4143), .C1(n196), .C2(n4178), .A(n1873), 
        .ZN(n1878) );
  OAI22_X1 U1525 ( .A1(n205), .A2(n1875), .B1(n202), .B2(n1874), .ZN(n1876) );
  AOI221_X1 U1526 ( .B1(n211), .B2(n4283), .C1(n208), .C2(n4341), .A(n1876), 
        .ZN(n1877) );
  NAND4_X1 U1527 ( .A1(n1880), .A2(n1879), .A3(n1878), .A4(n1877), .ZN(n1898)
         );
  OAI22_X1 U1528 ( .A1(n217), .A2(n1882), .B1(n214), .B2(n1881), .ZN(n1883) );
  AOI221_X1 U1529 ( .B1(n223), .B2(n2298), .C1(n220), .C2(n2332), .A(n1883), 
        .ZN(n1896) );
  OAI22_X1 U1530 ( .A1(n229), .A2(n1885), .B1(n226), .B2(n1884), .ZN(n1886) );
  AOI221_X1 U1531 ( .B1(n235), .B2(n2434), .C1(n232), .C2(n2472), .A(n1886), 
        .ZN(n1895) );
  OAI22_X1 U1532 ( .A1(n241), .A2(n1888), .B1(n238), .B2(n1887), .ZN(n1889) );
  AOI221_X1 U1533 ( .B1(n247), .B2(n2506), .C1(n244), .C2(n3628), .A(n1889), 
        .ZN(n1894) );
  OAI22_X1 U1534 ( .A1(n253), .A2(n1891), .B1(n250), .B2(n1890), .ZN(n1892) );
  AOI221_X1 U1535 ( .B1(n259), .B2(n3730), .C1(n256), .C2(n3764), .A(n1892), 
        .ZN(n1893) );
  NAND4_X1 U1536 ( .A1(n1896), .A2(n1895), .A3(n1894), .A4(n1893), .ZN(n1897)
         );
  OAI21_X1 U1537 ( .B1(n1898), .B2(n1897), .A(n262), .ZN(n1899) );
  OAI21_X1 U1538 ( .B1(n266), .B2(n1900), .A(n1899), .ZN(n2582) );
  OAI22_X1 U1539 ( .A1(n170), .A2(n1902), .B1(n167), .B2(n1901), .ZN(n1903) );
  AOI221_X1 U1540 ( .B1(n176), .B2(n3868), .C1(n173), .C2(n3902), .A(n1903), 
        .ZN(n1916) );
  OAI22_X1 U1541 ( .A1(n182), .A2(n1905), .B1(n179), .B2(n1904), .ZN(n1906) );
  AOI221_X1 U1542 ( .B1(n188), .B2(n4004), .C1(n185), .C2(n4038), .A(n1906), 
        .ZN(n1915) );
  OAI22_X1 U1543 ( .A1(n194), .A2(n1908), .B1(n191), .B2(n1907), .ZN(n1909) );
  AOI221_X1 U1544 ( .B1(n200), .B2(n4144), .C1(n197), .C2(n4179), .A(n1909), 
        .ZN(n1914) );
  OAI22_X1 U1545 ( .A1(n206), .A2(n1911), .B1(n203), .B2(n1910), .ZN(n1912) );
  AOI221_X1 U1546 ( .B1(n212), .B2(n4284), .C1(n209), .C2(n4343), .A(n1912), 
        .ZN(n1913) );
  NAND4_X1 U1547 ( .A1(n1916), .A2(n1915), .A3(n1914), .A4(n1913), .ZN(n1934)
         );
  OAI22_X1 U1548 ( .A1(n218), .A2(n1918), .B1(n215), .B2(n1917), .ZN(n1919) );
  AOI221_X1 U1549 ( .B1(n224), .B2(n2299), .C1(n221), .C2(n2333), .A(n1919), 
        .ZN(n1932) );
  OAI22_X1 U1550 ( .A1(n230), .A2(n1921), .B1(n227), .B2(n1920), .ZN(n1922) );
  AOI221_X1 U1551 ( .B1(n236), .B2(n2435), .C1(n233), .C2(n2473), .A(n1922), 
        .ZN(n1931) );
  OAI22_X1 U1552 ( .A1(n242), .A2(n1924), .B1(n239), .B2(n1923), .ZN(n1925) );
  AOI221_X1 U1553 ( .B1(n248), .B2(n2507), .C1(n245), .C2(n3629), .A(n1925), 
        .ZN(n1930) );
  OAI22_X1 U1554 ( .A1(n254), .A2(n1927), .B1(n251), .B2(n1926), .ZN(n1928) );
  AOI221_X1 U1555 ( .B1(n260), .B2(n3731), .C1(n257), .C2(n3765), .A(n1928), 
        .ZN(n1929) );
  NAND4_X1 U1556 ( .A1(n1932), .A2(n1931), .A3(n1930), .A4(n1929), .ZN(n1933)
         );
  OAI21_X1 U1557 ( .B1(n1934), .B2(n1933), .A(n263), .ZN(n1935) );
  OAI21_X1 U1558 ( .B1(n266), .B2(n1936), .A(n1935), .ZN(n2583) );
  OAI22_X1 U1559 ( .A1(n170), .A2(n1938), .B1(n167), .B2(n1937), .ZN(n1939) );
  AOI221_X1 U1560 ( .B1(n176), .B2(n3869), .C1(n173), .C2(n3903), .A(n1939), 
        .ZN(n1952) );
  OAI22_X1 U1561 ( .A1(n182), .A2(n1941), .B1(n179), .B2(n1940), .ZN(n1942) );
  AOI221_X1 U1562 ( .B1(n188), .B2(n4005), .C1(n185), .C2(n4039), .A(n1942), 
        .ZN(n1951) );
  OAI22_X1 U1563 ( .A1(n194), .A2(n1944), .B1(n191), .B2(n1943), .ZN(n1945) );
  AOI221_X1 U1564 ( .B1(n200), .B2(n4145), .C1(n197), .C2(n4180), .A(n1945), 
        .ZN(n1950) );
  OAI22_X1 U1565 ( .A1(n206), .A2(n1947), .B1(n203), .B2(n1946), .ZN(n1948) );
  AOI221_X1 U1566 ( .B1(n212), .B2(n4285), .C1(n209), .C2(n4345), .A(n1948), 
        .ZN(n1949) );
  NAND4_X1 U1567 ( .A1(n1952), .A2(n1951), .A3(n1950), .A4(n1949), .ZN(n1970)
         );
  OAI22_X1 U1568 ( .A1(n218), .A2(n1954), .B1(n215), .B2(n1953), .ZN(n1955) );
  AOI221_X1 U1569 ( .B1(n224), .B2(n2300), .C1(n221), .C2(n2334), .A(n1955), 
        .ZN(n1968) );
  OAI22_X1 U1570 ( .A1(n230), .A2(n1957), .B1(n227), .B2(n1956), .ZN(n1958) );
  AOI221_X1 U1571 ( .B1(n236), .B2(n2436), .C1(n233), .C2(n2474), .A(n1958), 
        .ZN(n1967) );
  OAI22_X1 U1572 ( .A1(n242), .A2(n1960), .B1(n239), .B2(n1959), .ZN(n1961) );
  AOI221_X1 U1573 ( .B1(n248), .B2(n2508), .C1(n245), .C2(n3630), .A(n1961), 
        .ZN(n1966) );
  OAI22_X1 U1574 ( .A1(n254), .A2(n1963), .B1(n251), .B2(n1962), .ZN(n1964) );
  AOI221_X1 U1575 ( .B1(n260), .B2(n3732), .C1(n257), .C2(n3766), .A(n1964), 
        .ZN(n1965) );
  NAND4_X1 U1576 ( .A1(n1968), .A2(n1967), .A3(n1966), .A4(n1965), .ZN(n1969)
         );
  OAI21_X1 U1577 ( .B1(n1970), .B2(n1969), .A(n263), .ZN(n1971) );
  OAI21_X1 U1578 ( .B1(n266), .B2(n1972), .A(n1971), .ZN(n2584) );
  OAI22_X1 U1579 ( .A1(n170), .A2(n1974), .B1(n167), .B2(n1973), .ZN(n1975) );
  AOI221_X1 U1580 ( .B1(n176), .B2(n3870), .C1(n173), .C2(n3904), .A(n1975), 
        .ZN(n1988) );
  OAI22_X1 U1581 ( .A1(n182), .A2(n1977), .B1(n179), .B2(n1976), .ZN(n1978) );
  AOI221_X1 U1582 ( .B1(n188), .B2(n4006), .C1(n185), .C2(n4040), .A(n1978), 
        .ZN(n1987) );
  OAI22_X1 U1583 ( .A1(n194), .A2(n1980), .B1(n191), .B2(n1979), .ZN(n1981) );
  AOI221_X1 U1584 ( .B1(n200), .B2(n4146), .C1(n197), .C2(n4181), .A(n1981), 
        .ZN(n1986) );
  OAI22_X1 U1585 ( .A1(n206), .A2(n1983), .B1(n203), .B2(n1982), .ZN(n1984) );
  AOI221_X1 U1586 ( .B1(n212), .B2(n4286), .C1(n209), .C2(n4347), .A(n1984), 
        .ZN(n1985) );
  NAND4_X1 U1587 ( .A1(n1988), .A2(n1987), .A3(n1986), .A4(n1985), .ZN(n2006)
         );
  OAI22_X1 U1588 ( .A1(n218), .A2(n1990), .B1(n215), .B2(n1989), .ZN(n1991) );
  AOI221_X1 U1589 ( .B1(n224), .B2(n2301), .C1(n221), .C2(n2335), .A(n1991), 
        .ZN(n2004) );
  OAI22_X1 U1590 ( .A1(n230), .A2(n1993), .B1(n227), .B2(n1992), .ZN(n1994) );
  AOI221_X1 U1591 ( .B1(n236), .B2(n2437), .C1(n233), .C2(n2475), .A(n1994), 
        .ZN(n2003) );
  OAI22_X1 U1592 ( .A1(n242), .A2(n1996), .B1(n239), .B2(n1995), .ZN(n1997) );
  AOI221_X1 U1593 ( .B1(n248), .B2(n2509), .C1(n245), .C2(n3631), .A(n1997), 
        .ZN(n2002) );
  OAI22_X1 U1594 ( .A1(n254), .A2(n1999), .B1(n251), .B2(n1998), .ZN(n2000) );
  AOI221_X1 U1595 ( .B1(n260), .B2(n3733), .C1(n257), .C2(n3767), .A(n2000), 
        .ZN(n2001) );
  NAND4_X1 U1596 ( .A1(n2004), .A2(n2003), .A3(n2002), .A4(n2001), .ZN(n2005)
         );
  OAI21_X1 U1597 ( .B1(n2006), .B2(n2005), .A(n263), .ZN(n2007) );
  OAI21_X1 U1598 ( .B1(n266), .B2(n2008), .A(n2007), .ZN(n2585) );
  OAI22_X1 U1599 ( .A1(n170), .A2(n2010), .B1(n167), .B2(n2009), .ZN(n2011) );
  AOI221_X1 U1600 ( .B1(n176), .B2(n3871), .C1(n173), .C2(n3905), .A(n2011), 
        .ZN(n2024) );
  OAI22_X1 U1601 ( .A1(n182), .A2(n2013), .B1(n179), .B2(n2012), .ZN(n2014) );
  AOI221_X1 U1602 ( .B1(n188), .B2(n4007), .C1(n185), .C2(n4041), .A(n2014), 
        .ZN(n2023) );
  OAI22_X1 U1603 ( .A1(n194), .A2(n2016), .B1(n191), .B2(n2015), .ZN(n2017) );
  AOI221_X1 U1604 ( .B1(n200), .B2(n4147), .C1(n197), .C2(n4182), .A(n2017), 
        .ZN(n2022) );
  OAI22_X1 U1605 ( .A1(n206), .A2(n2019), .B1(n203), .B2(n2018), .ZN(n2020) );
  AOI221_X1 U1606 ( .B1(n212), .B2(n4287), .C1(n209), .C2(n4349), .A(n2020), 
        .ZN(n2021) );
  NAND4_X1 U1607 ( .A1(n2024), .A2(n2023), .A3(n2022), .A4(n2021), .ZN(n2042)
         );
  OAI22_X1 U1608 ( .A1(n218), .A2(n2026), .B1(n215), .B2(n2025), .ZN(n2027) );
  AOI221_X1 U1609 ( .B1(n224), .B2(n2302), .C1(n221), .C2(n2336), .A(n2027), 
        .ZN(n2040) );
  OAI22_X1 U1610 ( .A1(n230), .A2(n2029), .B1(n227), .B2(n2028), .ZN(n2030) );
  AOI221_X1 U1611 ( .B1(n236), .B2(n2438), .C1(n233), .C2(n2476), .A(n2030), 
        .ZN(n2039) );
  OAI22_X1 U1612 ( .A1(n242), .A2(n2032), .B1(n239), .B2(n2031), .ZN(n2033) );
  AOI221_X1 U1613 ( .B1(n248), .B2(n2510), .C1(n245), .C2(n3632), .A(n2033), 
        .ZN(n2038) );
  OAI22_X1 U1614 ( .A1(n254), .A2(n2035), .B1(n251), .B2(n2034), .ZN(n2036) );
  AOI221_X1 U1615 ( .B1(n260), .B2(n3734), .C1(n257), .C2(n3768), .A(n2036), 
        .ZN(n2037) );
  NAND4_X1 U1616 ( .A1(n2040), .A2(n2039), .A3(n2038), .A4(n2037), .ZN(n2041)
         );
  OAI21_X1 U1617 ( .B1(n2042), .B2(n2041), .A(n263), .ZN(n2043) );
  OAI21_X1 U1618 ( .B1(n266), .B2(n2044), .A(n2043), .ZN(n2586) );
  OAI22_X1 U1619 ( .A1(n170), .A2(n2046), .B1(n167), .B2(n2045), .ZN(n2047) );
  AOI221_X1 U1620 ( .B1(n176), .B2(n3872), .C1(n173), .C2(n3906), .A(n2047), 
        .ZN(n2060) );
  OAI22_X1 U1621 ( .A1(n182), .A2(n2049), .B1(n179), .B2(n2048), .ZN(n2050) );
  AOI221_X1 U1622 ( .B1(n188), .B2(n4008), .C1(n185), .C2(n4042), .A(n2050), 
        .ZN(n2059) );
  OAI22_X1 U1623 ( .A1(n194), .A2(n2052), .B1(n191), .B2(n2051), .ZN(n2053) );
  AOI221_X1 U1624 ( .B1(n200), .B2(n4148), .C1(n197), .C2(n4183), .A(n2053), 
        .ZN(n2058) );
  OAI22_X1 U1625 ( .A1(n206), .A2(n2055), .B1(n203), .B2(n2054), .ZN(n2056) );
  AOI221_X1 U1626 ( .B1(n212), .B2(n4288), .C1(n209), .C2(n4351), .A(n2056), 
        .ZN(n2057) );
  NAND4_X1 U1627 ( .A1(n2060), .A2(n2059), .A3(n2058), .A4(n2057), .ZN(n2078)
         );
  OAI22_X1 U1628 ( .A1(n218), .A2(n2062), .B1(n215), .B2(n2061), .ZN(n2063) );
  AOI221_X1 U1629 ( .B1(n224), .B2(n2303), .C1(n221), .C2(n2337), .A(n2063), 
        .ZN(n2076) );
  OAI22_X1 U1630 ( .A1(n230), .A2(n2065), .B1(n227), .B2(n2064), .ZN(n2066) );
  AOI221_X1 U1631 ( .B1(n236), .B2(n2439), .C1(n233), .C2(n2477), .A(n2066), 
        .ZN(n2075) );
  OAI22_X1 U1632 ( .A1(n242), .A2(n2068), .B1(n239), .B2(n2067), .ZN(n2069) );
  AOI221_X1 U1633 ( .B1(n248), .B2(n2511), .C1(n245), .C2(n3633), .A(n2069), 
        .ZN(n2074) );
  OAI22_X1 U1634 ( .A1(n254), .A2(n2071), .B1(n251), .B2(n2070), .ZN(n2072) );
  AOI221_X1 U1635 ( .B1(n260), .B2(n3735), .C1(n257), .C2(n3769), .A(n2072), 
        .ZN(n2073) );
  NAND4_X1 U1636 ( .A1(n2076), .A2(n2075), .A3(n2074), .A4(n2073), .ZN(n2077)
         );
  OAI21_X1 U1637 ( .B1(n2078), .B2(n2077), .A(n263), .ZN(n2079) );
  OAI21_X1 U1638 ( .B1(n266), .B2(n2080), .A(n2079), .ZN(n2587) );
  OAI22_X1 U1639 ( .A1(n170), .A2(n2082), .B1(n167), .B2(n2081), .ZN(n2083) );
  AOI221_X1 U1640 ( .B1(n176), .B2(n3873), .C1(n173), .C2(n3907), .A(n2083), 
        .ZN(n2096) );
  OAI22_X1 U1641 ( .A1(n182), .A2(n2085), .B1(n179), .B2(n2084), .ZN(n2086) );
  AOI221_X1 U1642 ( .B1(n188), .B2(n4009), .C1(n185), .C2(n4043), .A(n2086), 
        .ZN(n2095) );
  OAI22_X1 U1643 ( .A1(n194), .A2(n2088), .B1(n191), .B2(n2087), .ZN(n2089) );
  AOI221_X1 U1644 ( .B1(n200), .B2(n4149), .C1(n197), .C2(n4184), .A(n2089), 
        .ZN(n2094) );
  OAI22_X1 U1645 ( .A1(n206), .A2(n2091), .B1(n203), .B2(n2090), .ZN(n2092) );
  AOI221_X1 U1646 ( .B1(n212), .B2(n4289), .C1(n209), .C2(n4353), .A(n2092), 
        .ZN(n2093) );
  NAND4_X1 U1647 ( .A1(n2096), .A2(n2095), .A3(n2094), .A4(n2093), .ZN(n2114)
         );
  OAI22_X1 U1648 ( .A1(n218), .A2(n2098), .B1(n215), .B2(n2097), .ZN(n2099) );
  AOI221_X1 U1649 ( .B1(n224), .B2(n2304), .C1(n221), .C2(n2338), .A(n2099), 
        .ZN(n2112) );
  OAI22_X1 U1650 ( .A1(n230), .A2(n2101), .B1(n227), .B2(n2100), .ZN(n2102) );
  AOI221_X1 U1651 ( .B1(n236), .B2(n2440), .C1(n233), .C2(n2478), .A(n2102), 
        .ZN(n2111) );
  OAI22_X1 U1652 ( .A1(n242), .A2(n2104), .B1(n239), .B2(n2103), .ZN(n2105) );
  AOI221_X1 U1653 ( .B1(n248), .B2(n2512), .C1(n245), .C2(n3634), .A(n2105), 
        .ZN(n2110) );
  OAI22_X1 U1654 ( .A1(n254), .A2(n2107), .B1(n251), .B2(n2106), .ZN(n2108) );
  AOI221_X1 U1655 ( .B1(n260), .B2(n3736), .C1(n257), .C2(n3770), .A(n2108), 
        .ZN(n2109) );
  NAND4_X1 U1656 ( .A1(n2112), .A2(n2111), .A3(n2110), .A4(n2109), .ZN(n2113)
         );
  OAI21_X1 U1657 ( .B1(n2114), .B2(n2113), .A(n263), .ZN(n2115) );
  OAI21_X1 U1658 ( .B1(n266), .B2(n2116), .A(n2115), .ZN(n2588) );
  OAI22_X1 U1659 ( .A1(n170), .A2(n2118), .B1(n167), .B2(n2117), .ZN(n2119) );
  AOI221_X1 U1660 ( .B1(n176), .B2(n3874), .C1(n173), .C2(n3908), .A(n2119), 
        .ZN(n2132) );
  OAI22_X1 U1661 ( .A1(n182), .A2(n2121), .B1(n179), .B2(n2120), .ZN(n2122) );
  AOI221_X1 U1662 ( .B1(n188), .B2(n4010), .C1(n185), .C2(n4044), .A(n2122), 
        .ZN(n2131) );
  OAI22_X1 U1663 ( .A1(n194), .A2(n2124), .B1(n191), .B2(n2123), .ZN(n2125) );
  AOI221_X1 U1664 ( .B1(n200), .B2(n4150), .C1(n197), .C2(n4185), .A(n2125), 
        .ZN(n2130) );
  OAI22_X1 U1665 ( .A1(n206), .A2(n2127), .B1(n203), .B2(n2126), .ZN(n2128) );
  AOI221_X1 U1666 ( .B1(n212), .B2(n4290), .C1(n209), .C2(n4355), .A(n2128), 
        .ZN(n2129) );
  NAND4_X1 U1667 ( .A1(n2132), .A2(n2131), .A3(n2130), .A4(n2129), .ZN(n2150)
         );
  OAI22_X1 U1668 ( .A1(n218), .A2(n2134), .B1(n215), .B2(n2133), .ZN(n2135) );
  AOI221_X1 U1669 ( .B1(n224), .B2(n2305), .C1(n221), .C2(n2339), .A(n2135), 
        .ZN(n2148) );
  OAI22_X1 U1670 ( .A1(n230), .A2(n2137), .B1(n227), .B2(n2136), .ZN(n2138) );
  AOI221_X1 U1671 ( .B1(n236), .B2(n2441), .C1(n233), .C2(n2479), .A(n2138), 
        .ZN(n2147) );
  OAI22_X1 U1672 ( .A1(n242), .A2(n2140), .B1(n239), .B2(n2139), .ZN(n2141) );
  AOI221_X1 U1673 ( .B1(n248), .B2(n2513), .C1(n245), .C2(n3635), .A(n2141), 
        .ZN(n2146) );
  OAI22_X1 U1674 ( .A1(n254), .A2(n2143), .B1(n251), .B2(n2142), .ZN(n2144) );
  AOI221_X1 U1675 ( .B1(n260), .B2(n3737), .C1(n257), .C2(n3771), .A(n2144), 
        .ZN(n2145) );
  NAND4_X1 U1676 ( .A1(n2148), .A2(n2147), .A3(n2146), .A4(n2145), .ZN(n2149)
         );
  OAI21_X1 U1677 ( .B1(n2150), .B2(n2149), .A(n263), .ZN(n2151) );
  OAI21_X1 U1678 ( .B1(n266), .B2(n2152), .A(n2151), .ZN(n2589) );
  OAI22_X1 U1679 ( .A1(n170), .A2(n2155), .B1(n167), .B2(n2153), .ZN(n2157) );
  AOI221_X1 U1680 ( .B1(n176), .B2(n3876), .C1(n173), .C2(n3910), .A(n2157), 
        .ZN(n2176) );
  OAI22_X1 U1681 ( .A1(n182), .A2(n2160), .B1(n179), .B2(n2158), .ZN(n2162) );
  AOI221_X1 U1682 ( .B1(n188), .B2(n4012), .C1(n185), .C2(n4046), .A(n2162), 
        .ZN(n2175) );
  OAI22_X1 U1683 ( .A1(n194), .A2(n2165), .B1(n191), .B2(n2163), .ZN(n2167) );
  AOI221_X1 U1684 ( .B1(n200), .B2(n4152), .C1(n197), .C2(n4187), .A(n2167), 
        .ZN(n2174) );
  OAI22_X1 U1685 ( .A1(n206), .A2(n2170), .B1(n203), .B2(n2168), .ZN(n2172) );
  AOI221_X1 U1686 ( .B1(n212), .B2(n4292), .C1(n209), .C2(n4358), .A(n2172), 
        .ZN(n2173) );
  NAND4_X1 U1687 ( .A1(n2176), .A2(n2175), .A3(n2174), .A4(n2173), .ZN(n2202)
         );
  OAI22_X1 U1688 ( .A1(n218), .A2(n2179), .B1(n215), .B2(n2177), .ZN(n2181) );
  AOI221_X1 U1689 ( .B1(n224), .B2(n2307), .C1(n221), .C2(n2341), .A(n2181), 
        .ZN(n2200) );
  OAI22_X1 U1690 ( .A1(n230), .A2(n2184), .B1(n227), .B2(n2182), .ZN(n2186) );
  AOI221_X1 U1691 ( .B1(n236), .B2(n2443), .C1(n233), .C2(n2481), .A(n2186), 
        .ZN(n2199) );
  OAI22_X1 U1692 ( .A1(n242), .A2(n2189), .B1(n239), .B2(n2187), .ZN(n2191) );
  AOI221_X1 U1693 ( .B1(n248), .B2(n2515), .C1(n245), .C2(n3637), .A(n2191), 
        .ZN(n2198) );
  OAI22_X1 U1694 ( .A1(n254), .A2(n2194), .B1(n251), .B2(n2192), .ZN(n2196) );
  AOI221_X1 U1695 ( .B1(n260), .B2(n3739), .C1(n257), .C2(n3773), .A(n2196), 
        .ZN(n2197) );
  NAND4_X1 U1696 ( .A1(n2200), .A2(n2199), .A3(n2198), .A4(n2197), .ZN(n2201)
         );
  OAI21_X1 U1697 ( .B1(n2202), .B2(n2201), .A(n263), .ZN(n2203) );
  OAI21_X1 U1698 ( .B1(n266), .B2(n2204), .A(n2203), .ZN(n2590) );
  NAND2_X1 U1699 ( .A1(DATAIN[0]), .A2(n368), .ZN(n4398) );
  NAND2_X1 U1700 ( .A1(n39), .A2(ADD_WR[0]), .ZN(n4118) );
  NAND2_X1 U1701 ( .A1(n62), .A2(ADD_WR[3]), .ZN(n2447) );
  OAI21_X1 U1702 ( .B1(n4118), .B2(n2447), .A(n363), .ZN(n2206) );
  INV_X1 U1703 ( .A(n2206), .ZN(n2238) );
  MUX2_X1 U1704 ( .A(n4398), .B(n1052), .S(n267), .Z(n2207) );
  INV_X1 U1705 ( .A(n2207), .ZN(n2591) );
  MUX2_X1 U1706 ( .A(n4400), .B(n1090), .S(n267), .Z(n2208) );
  INV_X1 U1707 ( .A(n2208), .ZN(n2592) );
  MUX2_X1 U1708 ( .A(n4402), .B(n1126), .S(n267), .Z(n2209) );
  INV_X1 U1709 ( .A(n2209), .ZN(n2593) );
  MUX2_X1 U1710 ( .A(n4404), .B(n1162), .S(n267), .Z(n2210) );
  INV_X1 U1711 ( .A(n2210), .ZN(n2594) );
  NAND2_X1 U1712 ( .A1(DATAIN[4]), .A2(n367), .ZN(n4406) );
  MUX2_X1 U1713 ( .A(n4406), .B(n1198), .S(n267), .Z(n2211) );
  INV_X1 U1714 ( .A(n2211), .ZN(n2595) );
  NAND2_X1 U1715 ( .A1(DATAIN[5]), .A2(n367), .ZN(n4408) );
  MUX2_X1 U1716 ( .A(n4408), .B(n1234), .S(n267), .Z(n2212) );
  INV_X1 U1717 ( .A(n2212), .ZN(n2596) );
  NAND2_X1 U1718 ( .A1(DATAIN[6]), .A2(n367), .ZN(n4410) );
  MUX2_X1 U1719 ( .A(n4410), .B(n1270), .S(n267), .Z(n2213) );
  INV_X1 U1720 ( .A(n2213), .ZN(n2597) );
  NAND2_X1 U1721 ( .A1(DATAIN[7]), .A2(n367), .ZN(n4412) );
  MUX2_X1 U1722 ( .A(n4412), .B(n1306), .S(n267), .Z(n2214) );
  INV_X1 U1723 ( .A(n2214), .ZN(n2598) );
  NAND2_X1 U1724 ( .A1(DATAIN[8]), .A2(n367), .ZN(n4414) );
  MUX2_X1 U1725 ( .A(n4414), .B(n1342), .S(n267), .Z(n2215) );
  INV_X1 U1726 ( .A(n2215), .ZN(n2599) );
  NAND2_X1 U1727 ( .A1(DATAIN[9]), .A2(n367), .ZN(n4416) );
  MUX2_X1 U1728 ( .A(n4416), .B(n1378), .S(n267), .Z(n2216) );
  INV_X1 U1729 ( .A(n2216), .ZN(n2600) );
  NAND2_X1 U1730 ( .A1(DATAIN[10]), .A2(n367), .ZN(n4418) );
  MUX2_X1 U1731 ( .A(n4418), .B(n1414), .S(n267), .Z(n2217) );
  INV_X1 U1732 ( .A(n2217), .ZN(n2601) );
  NAND2_X1 U1733 ( .A1(DATAIN[11]), .A2(n367), .ZN(n4420) );
  MUX2_X1 U1734 ( .A(n4420), .B(n1450), .S(n267), .Z(n2218) );
  INV_X1 U1735 ( .A(n2218), .ZN(n2602) );
  NAND2_X1 U1736 ( .A1(DATAIN[12]), .A2(n367), .ZN(n4422) );
  MUX2_X1 U1737 ( .A(n4422), .B(n1486), .S(n268), .Z(n2219) );
  INV_X1 U1738 ( .A(n2219), .ZN(n2603) );
  NAND2_X1 U1739 ( .A1(DATAIN[13]), .A2(n365), .ZN(n4424) );
  MUX2_X1 U1740 ( .A(n4424), .B(n1522), .S(n268), .Z(n2220) );
  INV_X1 U1741 ( .A(n2220), .ZN(n2604) );
  NAND2_X1 U1742 ( .A1(DATAIN[14]), .A2(n367), .ZN(n4426) );
  MUX2_X1 U1743 ( .A(n4426), .B(n1558), .S(n268), .Z(n2221) );
  INV_X1 U1744 ( .A(n2221), .ZN(n2605) );
  NAND2_X1 U1745 ( .A1(DATAIN[15]), .A2(n367), .ZN(n4428) );
  MUX2_X1 U1746 ( .A(n4428), .B(n1594), .S(n268), .Z(n2222) );
  INV_X1 U1747 ( .A(n2222), .ZN(n2606) );
  NAND2_X1 U1748 ( .A1(DATAIN[16]), .A2(n367), .ZN(n4430) );
  MUX2_X1 U1749 ( .A(n4430), .B(n1630), .S(n268), .Z(n2223) );
  INV_X1 U1750 ( .A(n2223), .ZN(n2607) );
  NAND2_X1 U1751 ( .A1(DATAIN[17]), .A2(n366), .ZN(n4432) );
  MUX2_X1 U1752 ( .A(n4432), .B(n1666), .S(n268), .Z(n2224) );
  INV_X1 U1753 ( .A(n2224), .ZN(n2608) );
  NAND2_X1 U1754 ( .A1(DATAIN[18]), .A2(n366), .ZN(n4434) );
  MUX2_X1 U1755 ( .A(n4434), .B(n1702), .S(n268), .Z(n2225) );
  INV_X1 U1756 ( .A(n2225), .ZN(n2609) );
  NAND2_X1 U1757 ( .A1(DATAIN[19]), .A2(n366), .ZN(n4436) );
  MUX2_X1 U1758 ( .A(n4436), .B(n1738), .S(n268), .Z(n2226) );
  INV_X1 U1759 ( .A(n2226), .ZN(n2610) );
  NAND2_X1 U1760 ( .A1(DATAIN[20]), .A2(n366), .ZN(n4438) );
  MUX2_X1 U1761 ( .A(n4438), .B(n1774), .S(n268), .Z(n2227) );
  INV_X1 U1762 ( .A(n2227), .ZN(n2611) );
  NAND2_X1 U1763 ( .A1(DATAIN[21]), .A2(n366), .ZN(n4440) );
  MUX2_X1 U1764 ( .A(n4440), .B(n1810), .S(n268), .Z(n2228) );
  INV_X1 U1765 ( .A(n2228), .ZN(n2612) );
  NAND2_X1 U1766 ( .A1(DATAIN[22]), .A2(n366), .ZN(n4442) );
  MUX2_X1 U1767 ( .A(n4442), .B(n1846), .S(n268), .Z(n2229) );
  INV_X1 U1768 ( .A(n2229), .ZN(n2613) );
  NAND2_X1 U1769 ( .A1(DATAIN[23]), .A2(n366), .ZN(n4444) );
  MUX2_X1 U1770 ( .A(n4444), .B(n1882), .S(n268), .Z(n2230) );
  INV_X1 U1771 ( .A(n2230), .ZN(n2614) );
  NAND2_X1 U1772 ( .A1(DATAIN[24]), .A2(n366), .ZN(n4446) );
  MUX2_X1 U1773 ( .A(n4446), .B(n1918), .S(n269), .Z(n2231) );
  INV_X1 U1774 ( .A(n2231), .ZN(n2615) );
  NAND2_X1 U1775 ( .A1(DATAIN[25]), .A2(n366), .ZN(n4448) );
  MUX2_X1 U1776 ( .A(n4448), .B(n1954), .S(n269), .Z(n2232) );
  INV_X1 U1777 ( .A(n2232), .ZN(n2616) );
  NAND2_X1 U1778 ( .A1(DATAIN[26]), .A2(n366), .ZN(n4450) );
  MUX2_X1 U1779 ( .A(n4450), .B(n1990), .S(n269), .Z(n2233) );
  INV_X1 U1780 ( .A(n2233), .ZN(n2617) );
  NAND2_X1 U1781 ( .A1(DATAIN[27]), .A2(n366), .ZN(n4452) );
  MUX2_X1 U1782 ( .A(n4452), .B(n2026), .S(n269), .Z(n2234) );
  INV_X1 U1783 ( .A(n2234), .ZN(n2618) );
  NAND2_X1 U1784 ( .A1(DATAIN[28]), .A2(n366), .ZN(n4454) );
  MUX2_X1 U1785 ( .A(n4454), .B(n2062), .S(n269), .Z(n2235) );
  INV_X1 U1786 ( .A(n2235), .ZN(n2619) );
  NAND2_X1 U1787 ( .A1(DATAIN[29]), .A2(n365), .ZN(n4456) );
  MUX2_X1 U1788 ( .A(n4456), .B(n2098), .S(n269), .Z(n2236) );
  INV_X1 U1789 ( .A(n2236), .ZN(n2620) );
  NAND2_X1 U1790 ( .A1(DATAIN[30]), .A2(n365), .ZN(n4458) );
  MUX2_X1 U1791 ( .A(n4458), .B(n2134), .S(n269), .Z(n2237) );
  INV_X1 U1792 ( .A(n2237), .ZN(n2621) );
  NAND2_X1 U1793 ( .A1(DATAIN[31]), .A2(n365), .ZN(n4461) );
  MUX2_X1 U1794 ( .A(n4461), .B(n2179), .S(n269), .Z(n2239) );
  INV_X1 U1795 ( .A(n2239), .ZN(n2622) );
  INV_X1 U1796 ( .A(ADD_WR[0]), .ZN(n2444) );
  NAND2_X1 U1797 ( .A1(n39), .A2(n2444), .ZN(n4153) );
  OAI21_X1 U1798 ( .B1(n4153), .B2(n2447), .A(n365), .ZN(n2240) );
  INV_X1 U1799 ( .A(n2240), .ZN(n2272) );
  MUX2_X1 U1800 ( .A(n4398), .B(n1051), .S(n270), .Z(n2241) );
  INV_X1 U1801 ( .A(n2241), .ZN(n2623) );
  MUX2_X1 U1802 ( .A(n4400), .B(n1089), .S(n270), .Z(n2242) );
  INV_X1 U1803 ( .A(n2242), .ZN(n2624) );
  MUX2_X1 U1804 ( .A(n4402), .B(n1125), .S(n270), .Z(n2243) );
  INV_X1 U1805 ( .A(n2243), .ZN(n2625) );
  MUX2_X1 U1806 ( .A(n4404), .B(n1161), .S(n270), .Z(n2244) );
  INV_X1 U1807 ( .A(n2244), .ZN(n2626) );
  MUX2_X1 U1808 ( .A(n4406), .B(n1197), .S(n270), .Z(n2245) );
  INV_X1 U1809 ( .A(n2245), .ZN(n2627) );
  MUX2_X1 U1810 ( .A(n4408), .B(n1233), .S(n270), .Z(n2246) );
  INV_X1 U1811 ( .A(n2246), .ZN(n2628) );
  MUX2_X1 U1812 ( .A(n4410), .B(n1269), .S(n270), .Z(n2247) );
  INV_X1 U1813 ( .A(n2247), .ZN(n2629) );
  MUX2_X1 U1814 ( .A(n4412), .B(n1305), .S(n270), .Z(n2248) );
  INV_X1 U1815 ( .A(n2248), .ZN(n2630) );
  MUX2_X1 U1816 ( .A(n4414), .B(n1341), .S(n270), .Z(n2249) );
  INV_X1 U1817 ( .A(n2249), .ZN(n2631) );
  MUX2_X1 U1818 ( .A(n4416), .B(n1377), .S(n270), .Z(n2250) );
  INV_X1 U1819 ( .A(n2250), .ZN(n2632) );
  MUX2_X1 U1820 ( .A(n4418), .B(n1413), .S(n270), .Z(n2251) );
  INV_X1 U1821 ( .A(n2251), .ZN(n2633) );
  MUX2_X1 U1822 ( .A(n4420), .B(n1449), .S(n270), .Z(n2252) );
  INV_X1 U1823 ( .A(n2252), .ZN(n2634) );
  MUX2_X1 U1824 ( .A(n4422), .B(n1485), .S(n271), .Z(n2253) );
  INV_X1 U1825 ( .A(n2253), .ZN(n2635) );
  MUX2_X1 U1826 ( .A(n4424), .B(n1521), .S(n271), .Z(n2254) );
  INV_X1 U1827 ( .A(n2254), .ZN(n2636) );
  MUX2_X1 U1828 ( .A(n4426), .B(n1557), .S(n271), .Z(n2255) );
  INV_X1 U1829 ( .A(n2255), .ZN(n2637) );
  MUX2_X1 U1830 ( .A(n4428), .B(n1593), .S(n271), .Z(n2256) );
  INV_X1 U1831 ( .A(n2256), .ZN(n2638) );
  MUX2_X1 U1832 ( .A(n4430), .B(n1629), .S(n271), .Z(n2257) );
  INV_X1 U1833 ( .A(n2257), .ZN(n2639) );
  MUX2_X1 U1834 ( .A(n4432), .B(n1665), .S(n271), .Z(n2258) );
  INV_X1 U1835 ( .A(n2258), .ZN(n2640) );
  MUX2_X1 U1836 ( .A(n4434), .B(n1701), .S(n271), .Z(n2259) );
  INV_X1 U1837 ( .A(n2259), .ZN(n2641) );
  MUX2_X1 U1838 ( .A(n4436), .B(n1737), .S(n271), .Z(n2260) );
  INV_X1 U1839 ( .A(n2260), .ZN(n2642) );
  MUX2_X1 U1840 ( .A(n4438), .B(n1773), .S(n271), .Z(n2261) );
  INV_X1 U1841 ( .A(n2261), .ZN(n2643) );
  MUX2_X1 U1842 ( .A(n4440), .B(n1809), .S(n271), .Z(n2262) );
  INV_X1 U1843 ( .A(n2262), .ZN(n2644) );
  MUX2_X1 U1844 ( .A(n4442), .B(n1845), .S(n271), .Z(n2263) );
  INV_X1 U1845 ( .A(n2263), .ZN(n2645) );
  MUX2_X1 U1846 ( .A(n4444), .B(n1881), .S(n271), .Z(n2264) );
  INV_X1 U1847 ( .A(n2264), .ZN(n2646) );
  MUX2_X1 U1848 ( .A(n4446), .B(n1917), .S(n272), .Z(n2265) );
  INV_X1 U1849 ( .A(n2265), .ZN(n2647) );
  MUX2_X1 U1850 ( .A(n4448), .B(n1953), .S(n272), .Z(n2266) );
  INV_X1 U1851 ( .A(n2266), .ZN(n2648) );
  MUX2_X1 U1852 ( .A(n4450), .B(n1989), .S(n272), .Z(n2267) );
  INV_X1 U1853 ( .A(n2267), .ZN(n2649) );
  MUX2_X1 U1854 ( .A(n4452), .B(n2025), .S(n272), .Z(n2268) );
  INV_X1 U1855 ( .A(n2268), .ZN(n2650) );
  MUX2_X1 U1856 ( .A(n4454), .B(n2061), .S(n272), .Z(n2269) );
  INV_X1 U1857 ( .A(n2269), .ZN(n2651) );
  MUX2_X1 U1858 ( .A(n4456), .B(n2097), .S(n272), .Z(n2270) );
  INV_X1 U1859 ( .A(n2270), .ZN(n2652) );
  MUX2_X1 U1860 ( .A(n4458), .B(n2133), .S(n272), .Z(n2271) );
  INV_X1 U1861 ( .A(n2271), .ZN(n2653) );
  MUX2_X1 U1862 ( .A(n4461), .B(n2177), .S(n272), .Z(n2273) );
  INV_X1 U1863 ( .A(n2273), .ZN(n2654) );
  INV_X1 U1864 ( .A(n4398), .ZN(n4296) );
  INV_X1 U1865 ( .A(ADD_WR[1]), .ZN(n2445) );
  NAND3_X1 U1866 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .A3(n2445), .ZN(n4188) );
  OAI21_X1 U1867 ( .B1(n4188), .B2(n2447), .A(n365), .ZN(n2274) );
  INV_X1 U1868 ( .A(n2274), .ZN(n2306) );
  MUX2_X1 U1869 ( .A(n4296), .B(n2275), .S(n273), .Z(n2655) );
  INV_X1 U1870 ( .A(n4400), .ZN(n4298) );
  MUX2_X1 U1871 ( .A(n4298), .B(n2276), .S(n273), .Z(n2656) );
  INV_X1 U1872 ( .A(n4402), .ZN(n4300) );
  MUX2_X1 U1873 ( .A(n4300), .B(n2277), .S(n273), .Z(n2657) );
  INV_X1 U1874 ( .A(n4404), .ZN(n4302) );
  MUX2_X1 U1875 ( .A(n4302), .B(n2278), .S(n273), .Z(n2658) );
  INV_X1 U1876 ( .A(n4406), .ZN(n4304) );
  MUX2_X1 U1877 ( .A(n4304), .B(n2279), .S(n273), .Z(n2659) );
  INV_X1 U1878 ( .A(n4408), .ZN(n4306) );
  MUX2_X1 U1879 ( .A(n4306), .B(n2280), .S(n273), .Z(n2660) );
  INV_X1 U1880 ( .A(n4410), .ZN(n4308) );
  MUX2_X1 U1881 ( .A(n4308), .B(n2281), .S(n273), .Z(n2661) );
  INV_X1 U1882 ( .A(n4412), .ZN(n4310) );
  MUX2_X1 U1883 ( .A(n4310), .B(n2282), .S(n273), .Z(n2662) );
  INV_X1 U1884 ( .A(n4414), .ZN(n4312) );
  MUX2_X1 U1885 ( .A(n4312), .B(n2283), .S(n273), .Z(n2663) );
  INV_X1 U1886 ( .A(n4416), .ZN(n4314) );
  MUX2_X1 U1887 ( .A(n4314), .B(n2284), .S(n273), .Z(n2664) );
  INV_X1 U1888 ( .A(n4418), .ZN(n4316) );
  MUX2_X1 U1889 ( .A(n4316), .B(n2285), .S(n273), .Z(n2665) );
  INV_X1 U1890 ( .A(n4420), .ZN(n4318) );
  MUX2_X1 U1891 ( .A(n4318), .B(n2286), .S(n273), .Z(n2666) );
  INV_X1 U1892 ( .A(n4422), .ZN(n4320) );
  MUX2_X1 U1893 ( .A(n4320), .B(n2287), .S(n274), .Z(n2667) );
  INV_X1 U1894 ( .A(n4424), .ZN(n4322) );
  MUX2_X1 U1895 ( .A(n4322), .B(n2288), .S(n274), .Z(n2668) );
  INV_X1 U1896 ( .A(n4426), .ZN(n4324) );
  MUX2_X1 U1897 ( .A(n4324), .B(n2289), .S(n274), .Z(n2669) );
  INV_X1 U1898 ( .A(n4428), .ZN(n4326) );
  MUX2_X1 U1899 ( .A(n4326), .B(n2290), .S(n274), .Z(n2670) );
  INV_X1 U1900 ( .A(n4430), .ZN(n4328) );
  MUX2_X1 U1901 ( .A(n4328), .B(n2291), .S(n274), .Z(n2671) );
  INV_X1 U1902 ( .A(n4432), .ZN(n4330) );
  MUX2_X1 U1903 ( .A(n4330), .B(n2292), .S(n274), .Z(n2672) );
  INV_X1 U1904 ( .A(n4434), .ZN(n4332) );
  MUX2_X1 U1905 ( .A(n4332), .B(n2293), .S(n274), .Z(n2673) );
  INV_X1 U1906 ( .A(n4436), .ZN(n4334) );
  MUX2_X1 U1907 ( .A(n4334), .B(n2294), .S(n274), .Z(n2674) );
  INV_X1 U1908 ( .A(n4438), .ZN(n4336) );
  MUX2_X1 U1909 ( .A(n4336), .B(n2295), .S(n274), .Z(n2675) );
  INV_X1 U1910 ( .A(n4440), .ZN(n4338) );
  MUX2_X1 U1911 ( .A(n4338), .B(n2296), .S(n274), .Z(n2676) );
  INV_X1 U1912 ( .A(n4442), .ZN(n4340) );
  MUX2_X1 U1913 ( .A(n4340), .B(n2297), .S(n274), .Z(n2677) );
  INV_X1 U1914 ( .A(n4444), .ZN(n4342) );
  MUX2_X1 U1915 ( .A(n4342), .B(n2298), .S(n274), .Z(n2678) );
  INV_X1 U1916 ( .A(n4446), .ZN(n4344) );
  MUX2_X1 U1917 ( .A(n4344), .B(n2299), .S(n275), .Z(n2679) );
  INV_X1 U1918 ( .A(n4448), .ZN(n4346) );
  MUX2_X1 U1919 ( .A(n4346), .B(n2300), .S(n275), .Z(n2680) );
  INV_X1 U1920 ( .A(n4450), .ZN(n4348) );
  MUX2_X1 U1921 ( .A(n4348), .B(n2301), .S(n275), .Z(n2681) );
  INV_X1 U1922 ( .A(n4452), .ZN(n4350) );
  MUX2_X1 U1923 ( .A(n4350), .B(n2302), .S(n275), .Z(n2682) );
  INV_X1 U1924 ( .A(n4454), .ZN(n4352) );
  MUX2_X1 U1925 ( .A(n4352), .B(n2303), .S(n275), .Z(n2683) );
  INV_X1 U1926 ( .A(n4456), .ZN(n4354) );
  MUX2_X1 U1927 ( .A(n4354), .B(n2304), .S(n275), .Z(n2684) );
  INV_X1 U1928 ( .A(n4458), .ZN(n4356) );
  MUX2_X1 U1929 ( .A(n4356), .B(n2305), .S(n275), .Z(n2685) );
  INV_X1 U1930 ( .A(n4461), .ZN(n4359) );
  MUX2_X1 U1931 ( .A(n4359), .B(n2307), .S(n275), .Z(n2686) );
  NAND3_X1 U1932 ( .A1(ADD_WR[2]), .A2(n2445), .A3(n2444), .ZN(n4223) );
  OAI21_X1 U1933 ( .B1(n4223), .B2(n2447), .A(n365), .ZN(n2308) );
  INV_X1 U1934 ( .A(n2308), .ZN(n2340) );
  MUX2_X1 U1935 ( .A(n4296), .B(n2309), .S(n276), .Z(n2687) );
  MUX2_X1 U1936 ( .A(n4298), .B(n2310), .S(n276), .Z(n2688) );
  MUX2_X1 U1937 ( .A(n4300), .B(n2311), .S(n276), .Z(n2689) );
  MUX2_X1 U1938 ( .A(n4302), .B(n2312), .S(n276), .Z(n2690) );
  MUX2_X1 U1939 ( .A(n4304), .B(n2313), .S(n276), .Z(n2691) );
  MUX2_X1 U1940 ( .A(n4306), .B(n2314), .S(n276), .Z(n2692) );
  MUX2_X1 U1941 ( .A(n4308), .B(n2315), .S(n276), .Z(n2693) );
  MUX2_X1 U1942 ( .A(n4310), .B(n2316), .S(n276), .Z(n2694) );
  MUX2_X1 U1943 ( .A(n4312), .B(n2317), .S(n276), .Z(n2695) );
  MUX2_X1 U1944 ( .A(n4314), .B(n2318), .S(n276), .Z(n2696) );
  MUX2_X1 U1945 ( .A(n4316), .B(n2319), .S(n276), .Z(n2697) );
  MUX2_X1 U1946 ( .A(n4318), .B(n2320), .S(n276), .Z(n2698) );
  MUX2_X1 U1947 ( .A(n4320), .B(n2321), .S(n277), .Z(n2699) );
  MUX2_X1 U1948 ( .A(n4322), .B(n2322), .S(n277), .Z(n2700) );
  MUX2_X1 U1949 ( .A(n4324), .B(n2323), .S(n277), .Z(n2701) );
  MUX2_X1 U1950 ( .A(n4326), .B(n2324), .S(n277), .Z(n2702) );
  MUX2_X1 U1951 ( .A(n4328), .B(n2325), .S(n277), .Z(n2703) );
  MUX2_X1 U1952 ( .A(n4330), .B(n2326), .S(n277), .Z(n2704) );
  MUX2_X1 U1953 ( .A(n4332), .B(n2327), .S(n277), .Z(n2705) );
  MUX2_X1 U1954 ( .A(n4334), .B(n2328), .S(n277), .Z(n2706) );
  MUX2_X1 U1955 ( .A(n4336), .B(n2329), .S(n277), .Z(n2707) );
  MUX2_X1 U1956 ( .A(n4338), .B(n2330), .S(n277), .Z(n2708) );
  MUX2_X1 U1957 ( .A(n4340), .B(n2331), .S(n277), .Z(n2709) );
  MUX2_X1 U1958 ( .A(n4342), .B(n2332), .S(n277), .Z(n2710) );
  MUX2_X1 U1959 ( .A(n4344), .B(n2333), .S(n278), .Z(n2711) );
  MUX2_X1 U1960 ( .A(n4346), .B(n2334), .S(n278), .Z(n2712) );
  MUX2_X1 U1961 ( .A(n4348), .B(n2335), .S(n278), .Z(n2713) );
  MUX2_X1 U1962 ( .A(n4350), .B(n2336), .S(n278), .Z(n2714) );
  MUX2_X1 U1963 ( .A(n4352), .B(n2337), .S(n278), .Z(n2715) );
  MUX2_X1 U1964 ( .A(n4354), .B(n2338), .S(n278), .Z(n2716) );
  MUX2_X1 U1965 ( .A(n4356), .B(n2339), .S(n278), .Z(n2717) );
  MUX2_X1 U1966 ( .A(n4359), .B(n2341), .S(n278), .Z(n2718) );
  INV_X1 U1967 ( .A(ADD_WR[2]), .ZN(n2446) );
  NAND3_X1 U1968 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(n2446), .ZN(n4258) );
  OAI21_X1 U1969 ( .B1(n4258), .B2(n2447), .A(n365), .ZN(n2342) );
  INV_X1 U1970 ( .A(n2342), .ZN(n2374) );
  MUX2_X1 U1971 ( .A(n4398), .B(n1055), .S(n279), .Z(n2343) );
  INV_X1 U1972 ( .A(n2343), .ZN(n2719) );
  MUX2_X1 U1973 ( .A(n4400), .B(n1093), .S(n279), .Z(n2344) );
  INV_X1 U1974 ( .A(n2344), .ZN(n2720) );
  MUX2_X1 U1975 ( .A(n4402), .B(n1129), .S(n279), .Z(n2345) );
  INV_X1 U1976 ( .A(n2345), .ZN(n2721) );
  MUX2_X1 U1977 ( .A(n4404), .B(n1165), .S(n279), .Z(n2346) );
  INV_X1 U1978 ( .A(n2346), .ZN(n2722) );
  MUX2_X1 U1979 ( .A(n4406), .B(n1201), .S(n279), .Z(n2347) );
  INV_X1 U1980 ( .A(n2347), .ZN(n2723) );
  MUX2_X1 U1981 ( .A(n4408), .B(n1237), .S(n279), .Z(n2348) );
  INV_X1 U1982 ( .A(n2348), .ZN(n2724) );
  MUX2_X1 U1983 ( .A(n4410), .B(n1273), .S(n279), .Z(n2349) );
  INV_X1 U1984 ( .A(n2349), .ZN(n2725) );
  MUX2_X1 U1985 ( .A(n4412), .B(n1309), .S(n279), .Z(n2350) );
  INV_X1 U1986 ( .A(n2350), .ZN(n2726) );
  MUX2_X1 U1987 ( .A(n4414), .B(n1345), .S(n279), .Z(n2351) );
  INV_X1 U1988 ( .A(n2351), .ZN(n2727) );
  MUX2_X1 U1989 ( .A(n4416), .B(n1381), .S(n279), .Z(n2352) );
  INV_X1 U1990 ( .A(n2352), .ZN(n2728) );
  MUX2_X1 U1991 ( .A(n4418), .B(n1417), .S(n279), .Z(n2353) );
  INV_X1 U1992 ( .A(n2353), .ZN(n2729) );
  MUX2_X1 U1993 ( .A(n4420), .B(n1453), .S(n279), .Z(n2354) );
  INV_X1 U1994 ( .A(n2354), .ZN(n2730) );
  MUX2_X1 U1995 ( .A(n4422), .B(n1489), .S(n280), .Z(n2355) );
  INV_X1 U1996 ( .A(n2355), .ZN(n2731) );
  MUX2_X1 U1997 ( .A(n4424), .B(n1525), .S(n280), .Z(n2356) );
  INV_X1 U1998 ( .A(n2356), .ZN(n2732) );
  MUX2_X1 U1999 ( .A(n4426), .B(n1561), .S(n280), .Z(n2357) );
  INV_X1 U2000 ( .A(n2357), .ZN(n2733) );
  MUX2_X1 U2001 ( .A(n4428), .B(n1597), .S(n280), .Z(n2358) );
  INV_X1 U2002 ( .A(n2358), .ZN(n2734) );
  MUX2_X1 U2003 ( .A(n4430), .B(n1633), .S(n280), .Z(n2359) );
  INV_X1 U2004 ( .A(n2359), .ZN(n2735) );
  MUX2_X1 U2005 ( .A(n4432), .B(n1669), .S(n280), .Z(n2360) );
  INV_X1 U2006 ( .A(n2360), .ZN(n2736) );
  MUX2_X1 U2007 ( .A(n4434), .B(n1705), .S(n280), .Z(n2361) );
  INV_X1 U2008 ( .A(n2361), .ZN(n2737) );
  MUX2_X1 U2009 ( .A(n4436), .B(n1741), .S(n280), .Z(n2362) );
  INV_X1 U2010 ( .A(n2362), .ZN(n2738) );
  MUX2_X1 U2011 ( .A(n4438), .B(n1777), .S(n280), .Z(n2363) );
  INV_X1 U2012 ( .A(n2363), .ZN(n2739) );
  MUX2_X1 U2013 ( .A(n4440), .B(n1813), .S(n280), .Z(n2364) );
  INV_X1 U2014 ( .A(n2364), .ZN(n2740) );
  MUX2_X1 U2015 ( .A(n4442), .B(n1849), .S(n280), .Z(n2365) );
  INV_X1 U2016 ( .A(n2365), .ZN(n2741) );
  MUX2_X1 U2017 ( .A(n4444), .B(n1885), .S(n280), .Z(n2366) );
  INV_X1 U2018 ( .A(n2366), .ZN(n2742) );
  MUX2_X1 U2019 ( .A(n4446), .B(n1921), .S(n281), .Z(n2367) );
  INV_X1 U2020 ( .A(n2367), .ZN(n2743) );
  MUX2_X1 U2021 ( .A(n4448), .B(n1957), .S(n281), .Z(n2368) );
  INV_X1 U2022 ( .A(n2368), .ZN(n2744) );
  MUX2_X1 U2023 ( .A(n4450), .B(n1993), .S(n281), .Z(n2369) );
  INV_X1 U2024 ( .A(n2369), .ZN(n2745) );
  MUX2_X1 U2025 ( .A(n4452), .B(n2029), .S(n281), .Z(n2370) );
  INV_X1 U2026 ( .A(n2370), .ZN(n2746) );
  MUX2_X1 U2027 ( .A(n4454), .B(n2065), .S(n281), .Z(n2371) );
  INV_X1 U2028 ( .A(n2371), .ZN(n2747) );
  MUX2_X1 U2029 ( .A(n4456), .B(n2101), .S(n281), .Z(n2372) );
  INV_X1 U2030 ( .A(n2372), .ZN(n2748) );
  MUX2_X1 U2031 ( .A(n4458), .B(n2137), .S(n281), .Z(n2373) );
  INV_X1 U2032 ( .A(n2373), .ZN(n2749) );
  MUX2_X1 U2033 ( .A(n4461), .B(n2184), .S(n281), .Z(n2375) );
  INV_X1 U2034 ( .A(n2375), .ZN(n2750) );
  NAND3_X1 U2035 ( .A1(ADD_WR[1]), .A2(n2446), .A3(n2444), .ZN(n4293) );
  OAI21_X1 U2036 ( .B1(n4293), .B2(n2447), .A(n365), .ZN(n2376) );
  INV_X1 U2037 ( .A(n2376), .ZN(n2408) );
  MUX2_X1 U2038 ( .A(n4398), .B(n1054), .S(n282), .Z(n2377) );
  INV_X1 U2039 ( .A(n2377), .ZN(n2751) );
  MUX2_X1 U2040 ( .A(n4400), .B(n1092), .S(n282), .Z(n2378) );
  INV_X1 U2041 ( .A(n2378), .ZN(n2752) );
  MUX2_X1 U2042 ( .A(n4402), .B(n1128), .S(n282), .Z(n2379) );
  INV_X1 U2043 ( .A(n2379), .ZN(n2753) );
  MUX2_X1 U2044 ( .A(n4404), .B(n1164), .S(n282), .Z(n2380) );
  INV_X1 U2045 ( .A(n2380), .ZN(n2754) );
  MUX2_X1 U2046 ( .A(n4406), .B(n1200), .S(n282), .Z(n2381) );
  INV_X1 U2047 ( .A(n2381), .ZN(n2755) );
  MUX2_X1 U2048 ( .A(n4408), .B(n1236), .S(n282), .Z(n2382) );
  INV_X1 U2049 ( .A(n2382), .ZN(n2756) );
  MUX2_X1 U2050 ( .A(n4410), .B(n1272), .S(n282), .Z(n2383) );
  INV_X1 U2051 ( .A(n2383), .ZN(n2757) );
  MUX2_X1 U2052 ( .A(n4412), .B(n1308), .S(n282), .Z(n2384) );
  INV_X1 U2053 ( .A(n2384), .ZN(n2758) );
  MUX2_X1 U2054 ( .A(n4414), .B(n1344), .S(n282), .Z(n2385) );
  INV_X1 U2055 ( .A(n2385), .ZN(n2759) );
  MUX2_X1 U2056 ( .A(n4416), .B(n1380), .S(n282), .Z(n2386) );
  INV_X1 U2057 ( .A(n2386), .ZN(n2760) );
  MUX2_X1 U2058 ( .A(n4418), .B(n1416), .S(n282), .Z(n2387) );
  INV_X1 U2059 ( .A(n2387), .ZN(n2761) );
  MUX2_X1 U2060 ( .A(n4420), .B(n1452), .S(n282), .Z(n2388) );
  INV_X1 U2061 ( .A(n2388), .ZN(n2762) );
  MUX2_X1 U2062 ( .A(n4422), .B(n1488), .S(n283), .Z(n2389) );
  INV_X1 U2063 ( .A(n2389), .ZN(n2763) );
  MUX2_X1 U2064 ( .A(n4424), .B(n1524), .S(n283), .Z(n2390) );
  INV_X1 U2065 ( .A(n2390), .ZN(n2764) );
  MUX2_X1 U2066 ( .A(n4426), .B(n1560), .S(n283), .Z(n2391) );
  INV_X1 U2067 ( .A(n2391), .ZN(n2765) );
  MUX2_X1 U2068 ( .A(n4428), .B(n1596), .S(n283), .Z(n2392) );
  INV_X1 U2069 ( .A(n2392), .ZN(n2766) );
  MUX2_X1 U2070 ( .A(n4430), .B(n1632), .S(n283), .Z(n2393) );
  INV_X1 U2071 ( .A(n2393), .ZN(n2767) );
  MUX2_X1 U2072 ( .A(n4432), .B(n1668), .S(n283), .Z(n2394) );
  INV_X1 U2073 ( .A(n2394), .ZN(n2768) );
  MUX2_X1 U2074 ( .A(n4434), .B(n1704), .S(n283), .Z(n2395) );
  INV_X1 U2075 ( .A(n2395), .ZN(n2769) );
  MUX2_X1 U2076 ( .A(n4436), .B(n1740), .S(n283), .Z(n2396) );
  INV_X1 U2077 ( .A(n2396), .ZN(n2770) );
  MUX2_X1 U2078 ( .A(n4438), .B(n1776), .S(n283), .Z(n2397) );
  INV_X1 U2079 ( .A(n2397), .ZN(n2771) );
  MUX2_X1 U2080 ( .A(n4440), .B(n1812), .S(n283), .Z(n2398) );
  INV_X1 U2081 ( .A(n2398), .ZN(n2772) );
  MUX2_X1 U2082 ( .A(n4442), .B(n1848), .S(n283), .Z(n2399) );
  INV_X1 U2083 ( .A(n2399), .ZN(n2773) );
  MUX2_X1 U2084 ( .A(n4444), .B(n1884), .S(n283), .Z(n2400) );
  INV_X1 U2085 ( .A(n2400), .ZN(n2774) );
  MUX2_X1 U2086 ( .A(n4446), .B(n1920), .S(n284), .Z(n2401) );
  INV_X1 U2087 ( .A(n2401), .ZN(n2775) );
  MUX2_X1 U2088 ( .A(n4448), .B(n1956), .S(n284), .Z(n2402) );
  INV_X1 U2089 ( .A(n2402), .ZN(n2776) );
  MUX2_X1 U2090 ( .A(n4450), .B(n1992), .S(n284), .Z(n2403) );
  INV_X1 U2091 ( .A(n2403), .ZN(n2777) );
  MUX2_X1 U2092 ( .A(n4452), .B(n2028), .S(n284), .Z(n2404) );
  INV_X1 U2093 ( .A(n2404), .ZN(n2778) );
  MUX2_X1 U2094 ( .A(n4454), .B(n2064), .S(n284), .Z(n2405) );
  INV_X1 U2095 ( .A(n2405), .ZN(n2779) );
  MUX2_X1 U2096 ( .A(n4456), .B(n2100), .S(n284), .Z(n2406) );
  INV_X1 U2097 ( .A(n2406), .ZN(n2780) );
  MUX2_X1 U2098 ( .A(n4458), .B(n2136), .S(n284), .Z(n2407) );
  INV_X1 U2099 ( .A(n2407), .ZN(n2781) );
  MUX2_X1 U2100 ( .A(n4461), .B(n2182), .S(n284), .Z(n2409) );
  INV_X1 U2101 ( .A(n2409), .ZN(n2782) );
  NAND3_X1 U2102 ( .A1(ADD_WR[0]), .A2(n2446), .A3(n2445), .ZN(n4360) );
  OAI21_X1 U2103 ( .B1(n4360), .B2(n2447), .A(n365), .ZN(n2410) );
  INV_X1 U2104 ( .A(n2410), .ZN(n2442) );
  MUX2_X1 U2105 ( .A(n4296), .B(n2411), .S(n285), .Z(n2783) );
  MUX2_X1 U2106 ( .A(n4298), .B(n2412), .S(n285), .Z(n2784) );
  MUX2_X1 U2107 ( .A(n4300), .B(n2413), .S(n285), .Z(n2785) );
  MUX2_X1 U2108 ( .A(n4302), .B(n2414), .S(n285), .Z(n2786) );
  MUX2_X1 U2109 ( .A(n4304), .B(n2415), .S(n285), .Z(n2787) );
  MUX2_X1 U2110 ( .A(n4306), .B(n2416), .S(n285), .Z(n2788) );
  MUX2_X1 U2111 ( .A(n4308), .B(n2417), .S(n285), .Z(n2789) );
  MUX2_X1 U2112 ( .A(n4310), .B(n2418), .S(n285), .Z(n2790) );
  MUX2_X1 U2113 ( .A(n4312), .B(n2419), .S(n285), .Z(n2791) );
  MUX2_X1 U2114 ( .A(n4314), .B(n2420), .S(n285), .Z(n2792) );
  MUX2_X1 U2115 ( .A(n4316), .B(n2421), .S(n285), .Z(n2793) );
  MUX2_X1 U2116 ( .A(n4318), .B(n2422), .S(n285), .Z(n2794) );
  MUX2_X1 U2117 ( .A(n4320), .B(n2423), .S(n286), .Z(n2795) );
  MUX2_X1 U2118 ( .A(n4322), .B(n2424), .S(n286), .Z(n2796) );
  MUX2_X1 U2119 ( .A(n4324), .B(n2425), .S(n286), .Z(n2797) );
  MUX2_X1 U2120 ( .A(n4326), .B(n2426), .S(n286), .Z(n2798) );
  MUX2_X1 U2121 ( .A(n4328), .B(n2427), .S(n286), .Z(n2799) );
  MUX2_X1 U2122 ( .A(n4330), .B(n2428), .S(n286), .Z(n2800) );
  MUX2_X1 U2123 ( .A(n4332), .B(n2429), .S(n286), .Z(n2801) );
  MUX2_X1 U2124 ( .A(n4334), .B(n2430), .S(n286), .Z(n2802) );
  MUX2_X1 U2125 ( .A(n4336), .B(n2431), .S(n286), .Z(n2803) );
  MUX2_X1 U2126 ( .A(n4338), .B(n2432), .S(n286), .Z(n2804) );
  MUX2_X1 U2127 ( .A(n4340), .B(n2433), .S(n286), .Z(n2805) );
  MUX2_X1 U2128 ( .A(n4342), .B(n2434), .S(n286), .Z(n2806) );
  MUX2_X1 U2129 ( .A(n4344), .B(n2435), .S(n287), .Z(n2807) );
  MUX2_X1 U2130 ( .A(n4346), .B(n2436), .S(n287), .Z(n2808) );
  MUX2_X1 U2131 ( .A(n4348), .B(n2437), .S(n287), .Z(n2809) );
  MUX2_X1 U2132 ( .A(n4350), .B(n2438), .S(n287), .Z(n2810) );
  MUX2_X1 U2133 ( .A(n4352), .B(n2439), .S(n287), .Z(n2811) );
  MUX2_X1 U2134 ( .A(n4354), .B(n2440), .S(n287), .Z(n2812) );
  MUX2_X1 U2135 ( .A(n4356), .B(n2441), .S(n287), .Z(n2813) );
  MUX2_X1 U2136 ( .A(n4359), .B(n2443), .S(n287), .Z(n2814) );
  NAND3_X1 U2137 ( .A1(n2446), .A2(n2445), .A3(n2444), .ZN(n4395) );
  OAI21_X1 U2138 ( .B1(n4395), .B2(n2447), .A(n365), .ZN(n2448) );
  INV_X1 U2139 ( .A(n2448), .ZN(n2480) );
  MUX2_X1 U2140 ( .A(n4296), .B(n2449), .S(n288), .Z(n2815) );
  MUX2_X1 U2141 ( .A(n4298), .B(n2450), .S(n288), .Z(n2816) );
  MUX2_X1 U2142 ( .A(n4300), .B(n2451), .S(n288), .Z(n2817) );
  MUX2_X1 U2143 ( .A(n4302), .B(n2452), .S(n288), .Z(n2818) );
  MUX2_X1 U2144 ( .A(n4304), .B(n2453), .S(n288), .Z(n2819) );
  MUX2_X1 U2145 ( .A(n4306), .B(n2454), .S(n288), .Z(n2820) );
  MUX2_X1 U2146 ( .A(n4308), .B(n2455), .S(n288), .Z(n2821) );
  MUX2_X1 U2147 ( .A(n4310), .B(n2456), .S(n288), .Z(n2822) );
  MUX2_X1 U2148 ( .A(n4312), .B(n2457), .S(n288), .Z(n2823) );
  MUX2_X1 U2149 ( .A(n4314), .B(n2458), .S(n288), .Z(n2824) );
  MUX2_X1 U2150 ( .A(n4316), .B(n2459), .S(n288), .Z(n2825) );
  MUX2_X1 U2151 ( .A(n4318), .B(n2460), .S(n288), .Z(n2826) );
  MUX2_X1 U2152 ( .A(n4320), .B(n2461), .S(n289), .Z(n2827) );
  MUX2_X1 U2153 ( .A(n4322), .B(n2462), .S(n289), .Z(n2828) );
  MUX2_X1 U2154 ( .A(n4324), .B(n2463), .S(n289), .Z(n2829) );
  MUX2_X1 U2155 ( .A(n4326), .B(n2464), .S(n289), .Z(n2830) );
  MUX2_X1 U2156 ( .A(n4328), .B(n2465), .S(n289), .Z(n2831) );
  MUX2_X1 U2157 ( .A(n4330), .B(n2466), .S(n289), .Z(n2832) );
  MUX2_X1 U2158 ( .A(n4332), .B(n2467), .S(n289), .Z(n2833) );
  MUX2_X1 U2159 ( .A(n4334), .B(n2468), .S(n289), .Z(n2834) );
  MUX2_X1 U2160 ( .A(n4336), .B(n2469), .S(n289), .Z(n2835) );
  MUX2_X1 U2161 ( .A(n4338), .B(n2470), .S(n289), .Z(n2836) );
  MUX2_X1 U2162 ( .A(n4340), .B(n2471), .S(n289), .Z(n2837) );
  MUX2_X1 U2163 ( .A(n4342), .B(n2472), .S(n289), .Z(n2838) );
  MUX2_X1 U2164 ( .A(n4344), .B(n2473), .S(n290), .Z(n2839) );
  MUX2_X1 U2165 ( .A(n4346), .B(n2474), .S(n290), .Z(n2840) );
  MUX2_X1 U2166 ( .A(n4348), .B(n2475), .S(n290), .Z(n2841) );
  MUX2_X1 U2167 ( .A(n4350), .B(n2476), .S(n290), .Z(n2842) );
  MUX2_X1 U2168 ( .A(n4352), .B(n2477), .S(n290), .Z(n2843) );
  MUX2_X1 U2169 ( .A(n4354), .B(n2478), .S(n290), .Z(n2844) );
  MUX2_X1 U2170 ( .A(n4356), .B(n2479), .S(n290), .Z(n2845) );
  MUX2_X1 U2171 ( .A(n4359), .B(n2481), .S(n290), .Z(n2846) );
  INV_X1 U2172 ( .A(ADD_WR[3]), .ZN(n4117) );
  NAND2_X1 U2173 ( .A1(n62), .A2(n4117), .ZN(n3808) );
  OAI21_X1 U2174 ( .B1(n4118), .B2(n3808), .A(n365), .ZN(n2482) );
  INV_X1 U2175 ( .A(n2482), .ZN(n2514) );
  MUX2_X1 U2176 ( .A(n4296), .B(n2483), .S(n291), .Z(n2847) );
  MUX2_X1 U2177 ( .A(n4298), .B(n2484), .S(n291), .Z(n2848) );
  MUX2_X1 U2178 ( .A(n4300), .B(n2485), .S(n291), .Z(n2849) );
  MUX2_X1 U2179 ( .A(n4302), .B(n2486), .S(n291), .Z(n2850) );
  MUX2_X1 U2180 ( .A(n4304), .B(n2487), .S(n291), .Z(n2851) );
  MUX2_X1 U2181 ( .A(n4306), .B(n2488), .S(n291), .Z(n2852) );
  MUX2_X1 U2182 ( .A(n4308), .B(n2489), .S(n291), .Z(n2853) );
  MUX2_X1 U2183 ( .A(n4310), .B(n2490), .S(n291), .Z(n2854) );
  MUX2_X1 U2184 ( .A(n4312), .B(n2491), .S(n291), .Z(n2855) );
  MUX2_X1 U2185 ( .A(n4314), .B(n2492), .S(n291), .Z(n2856) );
  MUX2_X1 U2186 ( .A(n4316), .B(n2493), .S(n291), .Z(n2857) );
  MUX2_X1 U2187 ( .A(n4318), .B(n2494), .S(n291), .Z(n2858) );
  MUX2_X1 U2188 ( .A(n4320), .B(n2495), .S(n292), .Z(n2859) );
  MUX2_X1 U2189 ( .A(n4322), .B(n2496), .S(n292), .Z(n2860) );
  MUX2_X1 U2190 ( .A(n4324), .B(n2497), .S(n292), .Z(n2861) );
  MUX2_X1 U2191 ( .A(n4326), .B(n2498), .S(n292), .Z(n2862) );
  MUX2_X1 U2192 ( .A(n4328), .B(n2499), .S(n292), .Z(n2863) );
  MUX2_X1 U2193 ( .A(n4330), .B(n2500), .S(n292), .Z(n2864) );
  MUX2_X1 U2194 ( .A(n4332), .B(n2501), .S(n292), .Z(n2865) );
  MUX2_X1 U2195 ( .A(n4334), .B(n2502), .S(n292), .Z(n2866) );
  MUX2_X1 U2196 ( .A(n4336), .B(n2503), .S(n292), .Z(n2867) );
  MUX2_X1 U2197 ( .A(n4338), .B(n2504), .S(n292), .Z(n2868) );
  MUX2_X1 U2198 ( .A(n4340), .B(n2505), .S(n292), .Z(n2869) );
  MUX2_X1 U2199 ( .A(n4342), .B(n2506), .S(n292), .Z(n2870) );
  MUX2_X1 U2200 ( .A(n4344), .B(n2507), .S(n293), .Z(n2871) );
  MUX2_X1 U2201 ( .A(n4346), .B(n2508), .S(n293), .Z(n2872) );
  MUX2_X1 U2202 ( .A(n4348), .B(n2509), .S(n293), .Z(n2873) );
  MUX2_X1 U2203 ( .A(n4350), .B(n2510), .S(n293), .Z(n2874) );
  MUX2_X1 U2204 ( .A(n4352), .B(n2511), .S(n293), .Z(n2875) );
  MUX2_X1 U2205 ( .A(n4354), .B(n2512), .S(n293), .Z(n2876) );
  MUX2_X1 U2206 ( .A(n4356), .B(n2513), .S(n293), .Z(n2877) );
  MUX2_X1 U2207 ( .A(n4359), .B(n2515), .S(n293), .Z(n2878) );
  OAI21_X1 U2208 ( .B1(n4153), .B2(n3808), .A(n364), .ZN(n2516) );
  INV_X1 U2209 ( .A(n2516), .ZN(n3636) );
  MUX2_X1 U2210 ( .A(n4296), .B(n2517), .S(n294), .Z(n2879) );
  MUX2_X1 U2211 ( .A(n4298), .B(n2518), .S(n294), .Z(n2880) );
  MUX2_X1 U2212 ( .A(n4300), .B(n2519), .S(n294), .Z(n2881) );
  MUX2_X1 U2213 ( .A(n4302), .B(n2520), .S(n294), .Z(n2882) );
  MUX2_X1 U2214 ( .A(n4304), .B(n2521), .S(n294), .Z(n2883) );
  MUX2_X1 U2215 ( .A(n4306), .B(n2522), .S(n294), .Z(n2884) );
  MUX2_X1 U2216 ( .A(n4308), .B(n2523), .S(n294), .Z(n2885) );
  MUX2_X1 U2217 ( .A(n4310), .B(n2524), .S(n294), .Z(n2886) );
  MUX2_X1 U2218 ( .A(n4312), .B(n2525), .S(n294), .Z(n2887) );
  MUX2_X1 U2219 ( .A(n4314), .B(n2526), .S(n294), .Z(n2888) );
  MUX2_X1 U2220 ( .A(n4316), .B(n3615), .S(n294), .Z(n2889) );
  MUX2_X1 U2221 ( .A(n4318), .B(n3616), .S(n294), .Z(n2890) );
  MUX2_X1 U2222 ( .A(n4320), .B(n3617), .S(n295), .Z(n2891) );
  MUX2_X1 U2223 ( .A(n4322), .B(n3618), .S(n295), .Z(n2892) );
  MUX2_X1 U2224 ( .A(n4324), .B(n3619), .S(n295), .Z(n2893) );
  MUX2_X1 U2225 ( .A(n4326), .B(n3620), .S(n295), .Z(n2894) );
  MUX2_X1 U2226 ( .A(n4328), .B(n3621), .S(n295), .Z(n2895) );
  MUX2_X1 U2227 ( .A(n4330), .B(n3622), .S(n295), .Z(n2896) );
  MUX2_X1 U2228 ( .A(n4332), .B(n3623), .S(n295), .Z(n2897) );
  MUX2_X1 U2229 ( .A(n4334), .B(n3624), .S(n295), .Z(n2898) );
  MUX2_X1 U2230 ( .A(n4336), .B(n3625), .S(n295), .Z(n2899) );
  MUX2_X1 U2231 ( .A(n4338), .B(n3626), .S(n295), .Z(n2900) );
  MUX2_X1 U2232 ( .A(n4340), .B(n3627), .S(n295), .Z(n2901) );
  MUX2_X1 U2233 ( .A(n4342), .B(n3628), .S(n295), .Z(n2902) );
  MUX2_X1 U2234 ( .A(n4344), .B(n3629), .S(n296), .Z(n2903) );
  MUX2_X1 U2235 ( .A(n4346), .B(n3630), .S(n296), .Z(n2904) );
  MUX2_X1 U2236 ( .A(n4348), .B(n3631), .S(n296), .Z(n2905) );
  MUX2_X1 U2237 ( .A(n4350), .B(n3632), .S(n296), .Z(n2906) );
  MUX2_X1 U2238 ( .A(n4352), .B(n3633), .S(n296), .Z(n2907) );
  MUX2_X1 U2239 ( .A(n4354), .B(n3634), .S(n296), .Z(n2908) );
  MUX2_X1 U2240 ( .A(n4356), .B(n3635), .S(n296), .Z(n2909) );
  MUX2_X1 U2241 ( .A(n4359), .B(n3637), .S(n296), .Z(n2910) );
  OAI21_X1 U2242 ( .B1(n4188), .B2(n3808), .A(n364), .ZN(n3638) );
  INV_X1 U2243 ( .A(n3638), .ZN(n3670) );
  MUX2_X1 U2244 ( .A(n4398), .B(n1060), .S(n297), .Z(n3639) );
  INV_X1 U2245 ( .A(n3639), .ZN(n2911) );
  MUX2_X1 U2246 ( .A(n4400), .B(n1096), .S(n297), .Z(n3640) );
  INV_X1 U2247 ( .A(n3640), .ZN(n2912) );
  MUX2_X1 U2248 ( .A(n4402), .B(n1132), .S(n297), .Z(n3641) );
  INV_X1 U2249 ( .A(n3641), .ZN(n2913) );
  MUX2_X1 U2250 ( .A(n4404), .B(n1168), .S(n297), .Z(n3642) );
  INV_X1 U2251 ( .A(n3642), .ZN(n2914) );
  MUX2_X1 U2252 ( .A(n4406), .B(n1204), .S(n297), .Z(n3643) );
  INV_X1 U2253 ( .A(n3643), .ZN(n2915) );
  MUX2_X1 U2254 ( .A(n4408), .B(n1240), .S(n297), .Z(n3644) );
  INV_X1 U2255 ( .A(n3644), .ZN(n2916) );
  MUX2_X1 U2256 ( .A(n4410), .B(n1276), .S(n297), .Z(n3645) );
  INV_X1 U2257 ( .A(n3645), .ZN(n2917) );
  MUX2_X1 U2258 ( .A(n4412), .B(n1312), .S(n297), .Z(n3646) );
  INV_X1 U2259 ( .A(n3646), .ZN(n2918) );
  MUX2_X1 U2260 ( .A(n4414), .B(n1348), .S(n297), .Z(n3647) );
  INV_X1 U2261 ( .A(n3647), .ZN(n2919) );
  MUX2_X1 U2262 ( .A(n4416), .B(n1384), .S(n297), .Z(n3648) );
  INV_X1 U2263 ( .A(n3648), .ZN(n2920) );
  MUX2_X1 U2264 ( .A(n4418), .B(n1420), .S(n297), .Z(n3649) );
  INV_X1 U2265 ( .A(n3649), .ZN(n2921) );
  MUX2_X1 U2266 ( .A(n4420), .B(n1456), .S(n297), .Z(n3650) );
  INV_X1 U2267 ( .A(n3650), .ZN(n2922) );
  MUX2_X1 U2268 ( .A(n4422), .B(n1492), .S(n298), .Z(n3651) );
  INV_X1 U2269 ( .A(n3651), .ZN(n2923) );
  MUX2_X1 U2270 ( .A(n4424), .B(n1528), .S(n298), .Z(n3652) );
  INV_X1 U2271 ( .A(n3652), .ZN(n2924) );
  MUX2_X1 U2272 ( .A(n4426), .B(n1564), .S(n298), .Z(n3653) );
  INV_X1 U2273 ( .A(n3653), .ZN(n2925) );
  MUX2_X1 U2274 ( .A(n4428), .B(n1600), .S(n298), .Z(n3654) );
  INV_X1 U2275 ( .A(n3654), .ZN(n2926) );
  MUX2_X1 U2276 ( .A(n4430), .B(n1636), .S(n298), .Z(n3655) );
  INV_X1 U2277 ( .A(n3655), .ZN(n2927) );
  MUX2_X1 U2278 ( .A(n4432), .B(n1672), .S(n298), .Z(n3656) );
  INV_X1 U2279 ( .A(n3656), .ZN(n2928) );
  MUX2_X1 U2280 ( .A(n4434), .B(n1708), .S(n298), .Z(n3657) );
  INV_X1 U2281 ( .A(n3657), .ZN(n2929) );
  MUX2_X1 U2282 ( .A(n4436), .B(n1744), .S(n298), .Z(n3658) );
  INV_X1 U2283 ( .A(n3658), .ZN(n2930) );
  MUX2_X1 U2284 ( .A(n4438), .B(n1780), .S(n298), .Z(n3659) );
  INV_X1 U2285 ( .A(n3659), .ZN(n2931) );
  MUX2_X1 U2286 ( .A(n4440), .B(n1816), .S(n298), .Z(n3660) );
  INV_X1 U2287 ( .A(n3660), .ZN(n2932) );
  MUX2_X1 U2288 ( .A(n4442), .B(n1852), .S(n298), .Z(n3661) );
  INV_X1 U2289 ( .A(n3661), .ZN(n2933) );
  MUX2_X1 U2290 ( .A(n4444), .B(n1888), .S(n298), .Z(n3662) );
  INV_X1 U2291 ( .A(n3662), .ZN(n2934) );
  MUX2_X1 U2292 ( .A(n4446), .B(n1924), .S(n299), .Z(n3663) );
  INV_X1 U2293 ( .A(n3663), .ZN(n2935) );
  MUX2_X1 U2294 ( .A(n4448), .B(n1960), .S(n299), .Z(n3664) );
  INV_X1 U2295 ( .A(n3664), .ZN(n2936) );
  MUX2_X1 U2296 ( .A(n4450), .B(n1996), .S(n299), .Z(n3665) );
  INV_X1 U2297 ( .A(n3665), .ZN(n2937) );
  MUX2_X1 U2298 ( .A(n4452), .B(n2032), .S(n299), .Z(n3666) );
  INV_X1 U2299 ( .A(n3666), .ZN(n2938) );
  MUX2_X1 U2300 ( .A(n4454), .B(n2068), .S(n299), .Z(n3667) );
  INV_X1 U2301 ( .A(n3667), .ZN(n2939) );
  MUX2_X1 U2302 ( .A(n4456), .B(n2104), .S(n299), .Z(n3668) );
  INV_X1 U2303 ( .A(n3668), .ZN(n2940) );
  MUX2_X1 U2304 ( .A(n4458), .B(n2140), .S(n299), .Z(n3669) );
  INV_X1 U2305 ( .A(n3669), .ZN(n2941) );
  MUX2_X1 U2306 ( .A(n4461), .B(n2189), .S(n299), .Z(n3671) );
  INV_X1 U2307 ( .A(n3671), .ZN(n2942) );
  OAI21_X1 U2308 ( .B1(n4223), .B2(n3808), .A(n364), .ZN(n3672) );
  INV_X1 U2309 ( .A(n3672), .ZN(n3704) );
  MUX2_X1 U2310 ( .A(n4398), .B(n1059), .S(n300), .Z(n3673) );
  INV_X1 U2311 ( .A(n3673), .ZN(n2943) );
  MUX2_X1 U2312 ( .A(n4400), .B(n1095), .S(n300), .Z(n3674) );
  INV_X1 U2313 ( .A(n3674), .ZN(n2944) );
  MUX2_X1 U2314 ( .A(n4402), .B(n1131), .S(n300), .Z(n3675) );
  INV_X1 U2315 ( .A(n3675), .ZN(n2945) );
  MUX2_X1 U2316 ( .A(n4404), .B(n1167), .S(n300), .Z(n3676) );
  INV_X1 U2317 ( .A(n3676), .ZN(n2946) );
  MUX2_X1 U2318 ( .A(n4406), .B(n1203), .S(n300), .Z(n3677) );
  INV_X1 U2319 ( .A(n3677), .ZN(n2947) );
  MUX2_X1 U2320 ( .A(n4408), .B(n1239), .S(n300), .Z(n3678) );
  INV_X1 U2321 ( .A(n3678), .ZN(n2948) );
  MUX2_X1 U2322 ( .A(n4410), .B(n1275), .S(n300), .Z(n3679) );
  INV_X1 U2323 ( .A(n3679), .ZN(n2949) );
  MUX2_X1 U2324 ( .A(n4412), .B(n1311), .S(n300), .Z(n3680) );
  INV_X1 U2325 ( .A(n3680), .ZN(n2950) );
  MUX2_X1 U2326 ( .A(n4414), .B(n1347), .S(n300), .Z(n3681) );
  INV_X1 U2327 ( .A(n3681), .ZN(n2951) );
  MUX2_X1 U2328 ( .A(n4416), .B(n1383), .S(n300), .Z(n3682) );
  INV_X1 U2329 ( .A(n3682), .ZN(n2952) );
  MUX2_X1 U2330 ( .A(n4418), .B(n1419), .S(n300), .Z(n3683) );
  INV_X1 U2331 ( .A(n3683), .ZN(n2953) );
  MUX2_X1 U2332 ( .A(n4420), .B(n1455), .S(n300), .Z(n3684) );
  INV_X1 U2333 ( .A(n3684), .ZN(n2954) );
  MUX2_X1 U2334 ( .A(n4422), .B(n1491), .S(n301), .Z(n3685) );
  INV_X1 U2335 ( .A(n3685), .ZN(n2955) );
  MUX2_X1 U2336 ( .A(n4424), .B(n1527), .S(n301), .Z(n3686) );
  INV_X1 U2337 ( .A(n3686), .ZN(n2956) );
  MUX2_X1 U2338 ( .A(n4426), .B(n1563), .S(n301), .Z(n3687) );
  INV_X1 U2339 ( .A(n3687), .ZN(n2957) );
  MUX2_X1 U2340 ( .A(n4428), .B(n1599), .S(n301), .Z(n3688) );
  INV_X1 U2341 ( .A(n3688), .ZN(n2958) );
  MUX2_X1 U2342 ( .A(n4430), .B(n1635), .S(n301), .Z(n3689) );
  INV_X1 U2343 ( .A(n3689), .ZN(n2959) );
  MUX2_X1 U2344 ( .A(n4432), .B(n1671), .S(n301), .Z(n3690) );
  INV_X1 U2345 ( .A(n3690), .ZN(n2960) );
  MUX2_X1 U2346 ( .A(n4434), .B(n1707), .S(n301), .Z(n3691) );
  INV_X1 U2347 ( .A(n3691), .ZN(n2961) );
  MUX2_X1 U2348 ( .A(n4436), .B(n1743), .S(n301), .Z(n3692) );
  INV_X1 U2349 ( .A(n3692), .ZN(n2962) );
  MUX2_X1 U2350 ( .A(n4438), .B(n1779), .S(n301), .Z(n3693) );
  INV_X1 U2351 ( .A(n3693), .ZN(n2963) );
  MUX2_X1 U2352 ( .A(n4440), .B(n1815), .S(n301), .Z(n3694) );
  INV_X1 U2353 ( .A(n3694), .ZN(n2964) );
  MUX2_X1 U2354 ( .A(n4442), .B(n1851), .S(n301), .Z(n3695) );
  INV_X1 U2355 ( .A(n3695), .ZN(n2965) );
  MUX2_X1 U2356 ( .A(n4444), .B(n1887), .S(n301), .Z(n3696) );
  INV_X1 U2357 ( .A(n3696), .ZN(n2966) );
  MUX2_X1 U2358 ( .A(n4446), .B(n1923), .S(n302), .Z(n3697) );
  INV_X1 U2359 ( .A(n3697), .ZN(n2967) );
  MUX2_X1 U2360 ( .A(n4448), .B(n1959), .S(n302), .Z(n3698) );
  INV_X1 U2361 ( .A(n3698), .ZN(n2968) );
  MUX2_X1 U2362 ( .A(n4450), .B(n1995), .S(n302), .Z(n3699) );
  INV_X1 U2363 ( .A(n3699), .ZN(n2969) );
  MUX2_X1 U2364 ( .A(n4452), .B(n2031), .S(n302), .Z(n3700) );
  INV_X1 U2365 ( .A(n3700), .ZN(n2970) );
  MUX2_X1 U2366 ( .A(n4454), .B(n2067), .S(n302), .Z(n3701) );
  INV_X1 U2367 ( .A(n3701), .ZN(n2971) );
  MUX2_X1 U2368 ( .A(n4456), .B(n2103), .S(n302), .Z(n3702) );
  INV_X1 U2369 ( .A(n3702), .ZN(n2972) );
  MUX2_X1 U2370 ( .A(n4458), .B(n2139), .S(n302), .Z(n3703) );
  INV_X1 U2371 ( .A(n3703), .ZN(n2973) );
  MUX2_X1 U2372 ( .A(n4461), .B(n2187), .S(n302), .Z(n3705) );
  INV_X1 U2373 ( .A(n3705), .ZN(n2974) );
  OAI21_X1 U2374 ( .B1(n4258), .B2(n3808), .A(n364), .ZN(n3706) );
  INV_X1 U2375 ( .A(n3706), .ZN(n3738) );
  MUX2_X1 U2376 ( .A(n4296), .B(n3707), .S(n303), .Z(n2975) );
  MUX2_X1 U2377 ( .A(n4298), .B(n3708), .S(n303), .Z(n2976) );
  MUX2_X1 U2378 ( .A(n4300), .B(n3709), .S(n303), .Z(n2977) );
  MUX2_X1 U2379 ( .A(n4302), .B(n3710), .S(n303), .Z(n2978) );
  MUX2_X1 U2380 ( .A(n4304), .B(n3711), .S(n303), .Z(n2979) );
  MUX2_X1 U2381 ( .A(n4306), .B(n3712), .S(n303), .Z(n2980) );
  MUX2_X1 U2382 ( .A(n4308), .B(n3713), .S(n303), .Z(n2981) );
  MUX2_X1 U2383 ( .A(n4310), .B(n3714), .S(n303), .Z(n2982) );
  MUX2_X1 U2384 ( .A(n4312), .B(n3715), .S(n303), .Z(n2983) );
  MUX2_X1 U2385 ( .A(n4314), .B(n3716), .S(n303), .Z(n2984) );
  MUX2_X1 U2386 ( .A(n4316), .B(n3717), .S(n303), .Z(n2985) );
  MUX2_X1 U2387 ( .A(n4318), .B(n3718), .S(n303), .Z(n2986) );
  MUX2_X1 U2388 ( .A(n4320), .B(n3719), .S(n304), .Z(n2987) );
  MUX2_X1 U2389 ( .A(n4322), .B(n3720), .S(n304), .Z(n2988) );
  MUX2_X1 U2390 ( .A(n4324), .B(n3721), .S(n304), .Z(n2989) );
  MUX2_X1 U2391 ( .A(n4326), .B(n3722), .S(n304), .Z(n2990) );
  MUX2_X1 U2392 ( .A(n4328), .B(n3723), .S(n304), .Z(n2991) );
  MUX2_X1 U2393 ( .A(n4330), .B(n3724), .S(n304), .Z(n2992) );
  MUX2_X1 U2394 ( .A(n4332), .B(n3725), .S(n304), .Z(n2993) );
  MUX2_X1 U2395 ( .A(n4334), .B(n3726), .S(n304), .Z(n2994) );
  MUX2_X1 U2396 ( .A(n4336), .B(n3727), .S(n304), .Z(n2995) );
  MUX2_X1 U2397 ( .A(n4338), .B(n3728), .S(n304), .Z(n2996) );
  MUX2_X1 U2398 ( .A(n4340), .B(n3729), .S(n304), .Z(n2997) );
  MUX2_X1 U2399 ( .A(n4342), .B(n3730), .S(n304), .Z(n2998) );
  MUX2_X1 U2400 ( .A(n4344), .B(n3731), .S(n305), .Z(n2999) );
  MUX2_X1 U2401 ( .A(n4346), .B(n3732), .S(n305), .Z(n3000) );
  MUX2_X1 U2402 ( .A(n4348), .B(n3733), .S(n305), .Z(n3001) );
  MUX2_X1 U2403 ( .A(n4350), .B(n3734), .S(n305), .Z(n3002) );
  MUX2_X1 U2404 ( .A(n4352), .B(n3735), .S(n305), .Z(n3003) );
  MUX2_X1 U2405 ( .A(n4354), .B(n3736), .S(n305), .Z(n3004) );
  MUX2_X1 U2406 ( .A(n4356), .B(n3737), .S(n305), .Z(n3005) );
  MUX2_X1 U2407 ( .A(n4359), .B(n3739), .S(n305), .Z(n3006) );
  OAI21_X1 U2408 ( .B1(n4293), .B2(n3808), .A(n364), .ZN(n3740) );
  INV_X1 U2409 ( .A(n3740), .ZN(n3772) );
  MUX2_X1 U2410 ( .A(n4296), .B(n3741), .S(n306), .Z(n3007) );
  MUX2_X1 U2411 ( .A(n4298), .B(n3742), .S(n306), .Z(n3008) );
  MUX2_X1 U2412 ( .A(n4300), .B(n3743), .S(n306), .Z(n3009) );
  MUX2_X1 U2413 ( .A(n4302), .B(n3744), .S(n306), .Z(n3010) );
  MUX2_X1 U2414 ( .A(n4304), .B(n3745), .S(n306), .Z(n3011) );
  MUX2_X1 U2415 ( .A(n4306), .B(n3746), .S(n306), .Z(n3012) );
  MUX2_X1 U2416 ( .A(n4308), .B(n3747), .S(n306), .Z(n3013) );
  MUX2_X1 U2417 ( .A(n4310), .B(n3748), .S(n306), .Z(n3014) );
  MUX2_X1 U2418 ( .A(n4312), .B(n3749), .S(n306), .Z(n3015) );
  MUX2_X1 U2419 ( .A(n4314), .B(n3750), .S(n306), .Z(n3016) );
  MUX2_X1 U2420 ( .A(n4316), .B(n3751), .S(n306), .Z(n3017) );
  MUX2_X1 U2421 ( .A(n4318), .B(n3752), .S(n306), .Z(n3018) );
  MUX2_X1 U2422 ( .A(n4320), .B(n3753), .S(n307), .Z(n3019) );
  MUX2_X1 U2423 ( .A(n4322), .B(n3754), .S(n307), .Z(n3020) );
  MUX2_X1 U2424 ( .A(n4324), .B(n3755), .S(n307), .Z(n3021) );
  MUX2_X1 U2425 ( .A(n4326), .B(n3756), .S(n307), .Z(n3022) );
  MUX2_X1 U2426 ( .A(n4328), .B(n3757), .S(n307), .Z(n3023) );
  MUX2_X1 U2427 ( .A(n4330), .B(n3758), .S(n307), .Z(n3024) );
  MUX2_X1 U2428 ( .A(n4332), .B(n3759), .S(n307), .Z(n3025) );
  MUX2_X1 U2429 ( .A(n4334), .B(n3760), .S(n307), .Z(n3026) );
  MUX2_X1 U2430 ( .A(n4336), .B(n3761), .S(n307), .Z(n3027) );
  MUX2_X1 U2431 ( .A(n4338), .B(n3762), .S(n307), .Z(n3028) );
  MUX2_X1 U2432 ( .A(n4340), .B(n3763), .S(n307), .Z(n3029) );
  MUX2_X1 U2433 ( .A(n4342), .B(n3764), .S(n307), .Z(n3030) );
  MUX2_X1 U2434 ( .A(n4344), .B(n3765), .S(n308), .Z(n3031) );
  MUX2_X1 U2435 ( .A(n4346), .B(n3766), .S(n308), .Z(n3032) );
  MUX2_X1 U2436 ( .A(n4348), .B(n3767), .S(n308), .Z(n3033) );
  MUX2_X1 U2437 ( .A(n4350), .B(n3768), .S(n308), .Z(n3034) );
  MUX2_X1 U2438 ( .A(n4352), .B(n3769), .S(n308), .Z(n3035) );
  MUX2_X1 U2439 ( .A(n4354), .B(n3770), .S(n308), .Z(n3036) );
  MUX2_X1 U2440 ( .A(n4356), .B(n3771), .S(n308), .Z(n3037) );
  MUX2_X1 U2441 ( .A(n4359), .B(n3773), .S(n308), .Z(n3038) );
  OAI21_X1 U2442 ( .B1(n4360), .B2(n3808), .A(n364), .ZN(n3774) );
  INV_X1 U2443 ( .A(n3774), .ZN(n3806) );
  MUX2_X1 U2444 ( .A(n4398), .B(n1063), .S(n309), .Z(n3775) );
  INV_X1 U2445 ( .A(n3775), .ZN(n3039) );
  MUX2_X1 U2446 ( .A(n4400), .B(n1099), .S(n309), .Z(n3776) );
  INV_X1 U2447 ( .A(n3776), .ZN(n3040) );
  MUX2_X1 U2448 ( .A(n4402), .B(n1135), .S(n309), .Z(n3777) );
  INV_X1 U2449 ( .A(n3777), .ZN(n3041) );
  MUX2_X1 U2450 ( .A(n4404), .B(n1171), .S(n309), .Z(n3778) );
  INV_X1 U2451 ( .A(n3778), .ZN(n3042) );
  MUX2_X1 U2452 ( .A(n4406), .B(n1207), .S(n309), .Z(n3779) );
  INV_X1 U2453 ( .A(n3779), .ZN(n3043) );
  MUX2_X1 U2454 ( .A(n4408), .B(n1243), .S(n309), .Z(n3780) );
  INV_X1 U2455 ( .A(n3780), .ZN(n3044) );
  MUX2_X1 U2456 ( .A(n4410), .B(n1279), .S(n309), .Z(n3781) );
  INV_X1 U2457 ( .A(n3781), .ZN(n3045) );
  MUX2_X1 U2458 ( .A(n4412), .B(n1315), .S(n309), .Z(n3782) );
  INV_X1 U2459 ( .A(n3782), .ZN(n3046) );
  MUX2_X1 U2460 ( .A(n4414), .B(n1351), .S(n309), .Z(n3783) );
  INV_X1 U2461 ( .A(n3783), .ZN(n3047) );
  MUX2_X1 U2462 ( .A(n4416), .B(n1387), .S(n309), .Z(n3784) );
  INV_X1 U2463 ( .A(n3784), .ZN(n3048) );
  MUX2_X1 U2464 ( .A(n4418), .B(n1423), .S(n309), .Z(n3785) );
  INV_X1 U2465 ( .A(n3785), .ZN(n3049) );
  MUX2_X1 U2466 ( .A(n4420), .B(n1459), .S(n309), .Z(n3786) );
  INV_X1 U2467 ( .A(n3786), .ZN(n3050) );
  MUX2_X1 U2468 ( .A(n4422), .B(n1495), .S(n310), .Z(n3787) );
  INV_X1 U2469 ( .A(n3787), .ZN(n3051) );
  MUX2_X1 U2470 ( .A(n4424), .B(n1531), .S(n310), .Z(n3788) );
  INV_X1 U2471 ( .A(n3788), .ZN(n3052) );
  MUX2_X1 U2472 ( .A(n4426), .B(n1567), .S(n310), .Z(n3789) );
  INV_X1 U2473 ( .A(n3789), .ZN(n3053) );
  MUX2_X1 U2474 ( .A(n4428), .B(n1603), .S(n310), .Z(n3790) );
  INV_X1 U2475 ( .A(n3790), .ZN(n3054) );
  MUX2_X1 U2476 ( .A(n4430), .B(n1639), .S(n310), .Z(n3791) );
  INV_X1 U2477 ( .A(n3791), .ZN(n3055) );
  MUX2_X1 U2478 ( .A(n4432), .B(n1675), .S(n310), .Z(n3792) );
  INV_X1 U2479 ( .A(n3792), .ZN(n3056) );
  MUX2_X1 U2480 ( .A(n4434), .B(n1711), .S(n310), .Z(n3793) );
  INV_X1 U2481 ( .A(n3793), .ZN(n3057) );
  MUX2_X1 U2482 ( .A(n4436), .B(n1747), .S(n310), .Z(n3794) );
  INV_X1 U2483 ( .A(n3794), .ZN(n3058) );
  MUX2_X1 U2484 ( .A(n4438), .B(n1783), .S(n310), .Z(n3795) );
  INV_X1 U2485 ( .A(n3795), .ZN(n3059) );
  MUX2_X1 U2486 ( .A(n4440), .B(n1819), .S(n310), .Z(n3796) );
  INV_X1 U2487 ( .A(n3796), .ZN(n3060) );
  MUX2_X1 U2488 ( .A(n4442), .B(n1855), .S(n310), .Z(n3797) );
  INV_X1 U2489 ( .A(n3797), .ZN(n3061) );
  MUX2_X1 U2490 ( .A(n4444), .B(n1891), .S(n310), .Z(n3798) );
  INV_X1 U2491 ( .A(n3798), .ZN(n3062) );
  MUX2_X1 U2492 ( .A(n4446), .B(n1927), .S(n311), .Z(n3799) );
  INV_X1 U2493 ( .A(n3799), .ZN(n3063) );
  MUX2_X1 U2494 ( .A(n4448), .B(n1963), .S(n311), .Z(n3800) );
  INV_X1 U2495 ( .A(n3800), .ZN(n3064) );
  MUX2_X1 U2496 ( .A(n4450), .B(n1999), .S(n311), .Z(n3801) );
  INV_X1 U2497 ( .A(n3801), .ZN(n3065) );
  MUX2_X1 U2498 ( .A(n4452), .B(n2035), .S(n311), .Z(n3802) );
  INV_X1 U2499 ( .A(n3802), .ZN(n3066) );
  MUX2_X1 U2500 ( .A(n4454), .B(n2071), .S(n311), .Z(n3803) );
  INV_X1 U2501 ( .A(n3803), .ZN(n3067) );
  MUX2_X1 U2502 ( .A(n4456), .B(n2107), .S(n311), .Z(n3804) );
  INV_X1 U2503 ( .A(n3804), .ZN(n3068) );
  MUX2_X1 U2504 ( .A(n4458), .B(n2143), .S(n311), .Z(n3805) );
  INV_X1 U2505 ( .A(n3805), .ZN(n3069) );
  MUX2_X1 U2506 ( .A(n4461), .B(n2194), .S(n311), .Z(n3807) );
  INV_X1 U2507 ( .A(n3807), .ZN(n3070) );
  OAI21_X1 U2508 ( .B1(n4395), .B2(n3808), .A(n364), .ZN(n3809) );
  INV_X1 U2509 ( .A(n3809), .ZN(n3841) );
  MUX2_X1 U2510 ( .A(n4398), .B(n1062), .S(n312), .Z(n3810) );
  INV_X1 U2511 ( .A(n3810), .ZN(n3071) );
  MUX2_X1 U2512 ( .A(n4400), .B(n1098), .S(n312), .Z(n3811) );
  INV_X1 U2513 ( .A(n3811), .ZN(n3072) );
  MUX2_X1 U2514 ( .A(n4402), .B(n1134), .S(n312), .Z(n3812) );
  INV_X1 U2515 ( .A(n3812), .ZN(n3073) );
  MUX2_X1 U2516 ( .A(n4404), .B(n1170), .S(n312), .Z(n3813) );
  INV_X1 U2517 ( .A(n3813), .ZN(n3074) );
  MUX2_X1 U2518 ( .A(n4406), .B(n1206), .S(n312), .Z(n3814) );
  INV_X1 U2519 ( .A(n3814), .ZN(n3075) );
  MUX2_X1 U2520 ( .A(n4408), .B(n1242), .S(n312), .Z(n3815) );
  INV_X1 U2521 ( .A(n3815), .ZN(n3076) );
  MUX2_X1 U2522 ( .A(n4410), .B(n1278), .S(n312), .Z(n3816) );
  INV_X1 U2523 ( .A(n3816), .ZN(n3077) );
  MUX2_X1 U2524 ( .A(n4412), .B(n1314), .S(n312), .Z(n3817) );
  INV_X1 U2525 ( .A(n3817), .ZN(n3078) );
  MUX2_X1 U2526 ( .A(n4414), .B(n1350), .S(n312), .Z(n3818) );
  INV_X1 U2527 ( .A(n3818), .ZN(n3079) );
  MUX2_X1 U2528 ( .A(n4416), .B(n1386), .S(n312), .Z(n3819) );
  INV_X1 U2529 ( .A(n3819), .ZN(n3080) );
  MUX2_X1 U2530 ( .A(n4418), .B(n1422), .S(n312), .Z(n3820) );
  INV_X1 U2531 ( .A(n3820), .ZN(n3081) );
  MUX2_X1 U2532 ( .A(n4420), .B(n1458), .S(n312), .Z(n3821) );
  INV_X1 U2533 ( .A(n3821), .ZN(n3082) );
  MUX2_X1 U2534 ( .A(n4422), .B(n1494), .S(n313), .Z(n3822) );
  INV_X1 U2535 ( .A(n3822), .ZN(n3083) );
  MUX2_X1 U2536 ( .A(n4424), .B(n1530), .S(n313), .Z(n3823) );
  INV_X1 U2537 ( .A(n3823), .ZN(n3084) );
  MUX2_X1 U2538 ( .A(n4426), .B(n1566), .S(n313), .Z(n3824) );
  INV_X1 U2539 ( .A(n3824), .ZN(n3085) );
  MUX2_X1 U2540 ( .A(n4428), .B(n1602), .S(n313), .Z(n3825) );
  INV_X1 U2541 ( .A(n3825), .ZN(n3086) );
  MUX2_X1 U2542 ( .A(n4430), .B(n1638), .S(n313), .Z(n3826) );
  INV_X1 U2543 ( .A(n3826), .ZN(n3087) );
  MUX2_X1 U2544 ( .A(n4432), .B(n1674), .S(n313), .Z(n3827) );
  INV_X1 U2545 ( .A(n3827), .ZN(n3088) );
  MUX2_X1 U2546 ( .A(n4434), .B(n1710), .S(n313), .Z(n3828) );
  INV_X1 U2547 ( .A(n3828), .ZN(n3089) );
  MUX2_X1 U2548 ( .A(n4436), .B(n1746), .S(n313), .Z(n3829) );
  INV_X1 U2549 ( .A(n3829), .ZN(n3090) );
  MUX2_X1 U2550 ( .A(n4438), .B(n1782), .S(n313), .Z(n3830) );
  INV_X1 U2551 ( .A(n3830), .ZN(n3091) );
  MUX2_X1 U2552 ( .A(n4440), .B(n1818), .S(n313), .Z(n3831) );
  INV_X1 U2553 ( .A(n3831), .ZN(n3092) );
  MUX2_X1 U2554 ( .A(n4442), .B(n1854), .S(n313), .Z(n3832) );
  INV_X1 U2555 ( .A(n3832), .ZN(n3093) );
  MUX2_X1 U2556 ( .A(n4444), .B(n1890), .S(n313), .Z(n3833) );
  INV_X1 U2557 ( .A(n3833), .ZN(n3094) );
  MUX2_X1 U2558 ( .A(n4446), .B(n1926), .S(n314), .Z(n3834) );
  INV_X1 U2559 ( .A(n3834), .ZN(n3095) );
  MUX2_X1 U2560 ( .A(n4448), .B(n1962), .S(n314), .Z(n3835) );
  INV_X1 U2561 ( .A(n3835), .ZN(n3096) );
  MUX2_X1 U2562 ( .A(n4450), .B(n1998), .S(n314), .Z(n3836) );
  INV_X1 U2563 ( .A(n3836), .ZN(n3097) );
  MUX2_X1 U2564 ( .A(n4452), .B(n2034), .S(n314), .Z(n3837) );
  INV_X1 U2565 ( .A(n3837), .ZN(n3098) );
  MUX2_X1 U2566 ( .A(n4454), .B(n2070), .S(n314), .Z(n3838) );
  INV_X1 U2567 ( .A(n3838), .ZN(n3099) );
  MUX2_X1 U2568 ( .A(n4456), .B(n2106), .S(n314), .Z(n3839) );
  INV_X1 U2569 ( .A(n3839), .ZN(n3100) );
  MUX2_X1 U2570 ( .A(n4458), .B(n2142), .S(n314), .Z(n3840) );
  INV_X1 U2571 ( .A(n3840), .ZN(n3101) );
  MUX2_X1 U2572 ( .A(n4461), .B(n2192), .S(n314), .Z(n3842) );
  INV_X1 U2573 ( .A(n3842), .ZN(n3102) );
  INV_X1 U2574 ( .A(ADD_WR[4]), .ZN(n4116) );
  NAND3_X1 U2575 ( .A1(ADD_WR[3]), .A2(WR), .A3(n4116), .ZN(n4081) );
  OAI21_X1 U2576 ( .B1(n4118), .B2(n4081), .A(n364), .ZN(n3843) );
  INV_X1 U2577 ( .A(n3843), .ZN(n3875) );
  MUX2_X1 U2578 ( .A(n4296), .B(n3844), .S(n315), .Z(n3103) );
  MUX2_X1 U2579 ( .A(n4298), .B(n3845), .S(n315), .Z(n3104) );
  MUX2_X1 U2580 ( .A(n4300), .B(n3846), .S(n315), .Z(n3105) );
  MUX2_X1 U2581 ( .A(n4302), .B(n3847), .S(n315), .Z(n3106) );
  MUX2_X1 U2582 ( .A(n4304), .B(n3848), .S(n315), .Z(n3107) );
  MUX2_X1 U2583 ( .A(n4306), .B(n3849), .S(n315), .Z(n3108) );
  MUX2_X1 U2584 ( .A(n4308), .B(n3850), .S(n315), .Z(n3109) );
  MUX2_X1 U2585 ( .A(n4310), .B(n3851), .S(n315), .Z(n3110) );
  MUX2_X1 U2586 ( .A(n4312), .B(n3852), .S(n315), .Z(n3111) );
  MUX2_X1 U2587 ( .A(n4314), .B(n3853), .S(n315), .Z(n3112) );
  MUX2_X1 U2588 ( .A(n4316), .B(n3854), .S(n315), .Z(n3113) );
  MUX2_X1 U2589 ( .A(n4318), .B(n3855), .S(n315), .Z(n3114) );
  MUX2_X1 U2590 ( .A(n4320), .B(n3856), .S(n316), .Z(n3115) );
  MUX2_X1 U2591 ( .A(n4322), .B(n3857), .S(n316), .Z(n3116) );
  MUX2_X1 U2592 ( .A(n4324), .B(n3858), .S(n316), .Z(n3117) );
  MUX2_X1 U2593 ( .A(n4326), .B(n3859), .S(n316), .Z(n3118) );
  MUX2_X1 U2594 ( .A(n4328), .B(n3860), .S(n316), .Z(n3119) );
  MUX2_X1 U2595 ( .A(n4330), .B(n3861), .S(n316), .Z(n3120) );
  MUX2_X1 U2596 ( .A(n4332), .B(n3862), .S(n316), .Z(n3121) );
  MUX2_X1 U2597 ( .A(n4334), .B(n3863), .S(n316), .Z(n3122) );
  MUX2_X1 U2598 ( .A(n4336), .B(n3864), .S(n316), .Z(n3123) );
  MUX2_X1 U2599 ( .A(n4338), .B(n3865), .S(n316), .Z(n3124) );
  MUX2_X1 U2600 ( .A(n4340), .B(n3866), .S(n316), .Z(n3125) );
  MUX2_X1 U2601 ( .A(n4342), .B(n3867), .S(n316), .Z(n3126) );
  MUX2_X1 U2602 ( .A(n4344), .B(n3868), .S(n317), .Z(n3127) );
  MUX2_X1 U2603 ( .A(n4346), .B(n3869), .S(n317), .Z(n3128) );
  MUX2_X1 U2604 ( .A(n4348), .B(n3870), .S(n317), .Z(n3129) );
  MUX2_X1 U2605 ( .A(n4350), .B(n3871), .S(n317), .Z(n3130) );
  MUX2_X1 U2606 ( .A(n4352), .B(n3872), .S(n317), .Z(n3131) );
  MUX2_X1 U2607 ( .A(n4354), .B(n3873), .S(n317), .Z(n3132) );
  MUX2_X1 U2608 ( .A(n4356), .B(n3874), .S(n317), .Z(n3133) );
  MUX2_X1 U2609 ( .A(n4359), .B(n3876), .S(n317), .Z(n3134) );
  OAI21_X1 U2610 ( .B1(n4153), .B2(n4081), .A(n364), .ZN(n3877) );
  INV_X1 U2611 ( .A(n3877), .ZN(n3909) );
  MUX2_X1 U2612 ( .A(n4296), .B(n3878), .S(n318), .Z(n3135) );
  MUX2_X1 U2613 ( .A(n4298), .B(n3879), .S(n318), .Z(n3136) );
  MUX2_X1 U2614 ( .A(n4300), .B(n3880), .S(n318), .Z(n3137) );
  MUX2_X1 U2615 ( .A(n4302), .B(n3881), .S(n318), .Z(n3138) );
  MUX2_X1 U2616 ( .A(n4304), .B(n3882), .S(n318), .Z(n3139) );
  MUX2_X1 U2617 ( .A(n4306), .B(n3883), .S(n318), .Z(n3140) );
  MUX2_X1 U2618 ( .A(n4308), .B(n3884), .S(n318), .Z(n3141) );
  MUX2_X1 U2619 ( .A(n4310), .B(n3885), .S(n318), .Z(n3142) );
  MUX2_X1 U2620 ( .A(n4312), .B(n3886), .S(n318), .Z(n3143) );
  MUX2_X1 U2621 ( .A(n4314), .B(n3887), .S(n318), .Z(n3144) );
  MUX2_X1 U2622 ( .A(n4316), .B(n3888), .S(n318), .Z(n3145) );
  MUX2_X1 U2623 ( .A(n4318), .B(n3889), .S(n318), .Z(n3146) );
  MUX2_X1 U2624 ( .A(n4320), .B(n3890), .S(n319), .Z(n3147) );
  MUX2_X1 U2625 ( .A(n4322), .B(n3891), .S(n319), .Z(n3148) );
  MUX2_X1 U2626 ( .A(n4324), .B(n3892), .S(n319), .Z(n3149) );
  MUX2_X1 U2627 ( .A(n4326), .B(n3893), .S(n319), .Z(n3150) );
  MUX2_X1 U2628 ( .A(n4328), .B(n3894), .S(n319), .Z(n3151) );
  MUX2_X1 U2629 ( .A(n4330), .B(n3895), .S(n319), .Z(n3152) );
  MUX2_X1 U2630 ( .A(n4332), .B(n3896), .S(n319), .Z(n3153) );
  MUX2_X1 U2631 ( .A(n4334), .B(n3897), .S(n319), .Z(n3154) );
  MUX2_X1 U2632 ( .A(n4336), .B(n3898), .S(n319), .Z(n3155) );
  MUX2_X1 U2633 ( .A(n4338), .B(n3899), .S(n319), .Z(n3156) );
  MUX2_X1 U2634 ( .A(n4340), .B(n3900), .S(n319), .Z(n3157) );
  MUX2_X1 U2635 ( .A(n4342), .B(n3901), .S(n319), .Z(n3158) );
  MUX2_X1 U2636 ( .A(n4344), .B(n3902), .S(n320), .Z(n3159) );
  MUX2_X1 U2637 ( .A(n4346), .B(n3903), .S(n320), .Z(n3160) );
  MUX2_X1 U2638 ( .A(n4348), .B(n3904), .S(n320), .Z(n3161) );
  MUX2_X1 U2639 ( .A(n4350), .B(n3905), .S(n320), .Z(n3162) );
  MUX2_X1 U2640 ( .A(n4352), .B(n3906), .S(n320), .Z(n3163) );
  MUX2_X1 U2641 ( .A(n4354), .B(n3907), .S(n320), .Z(n3164) );
  MUX2_X1 U2642 ( .A(n4356), .B(n3908), .S(n320), .Z(n3165) );
  MUX2_X1 U2643 ( .A(n4359), .B(n3910), .S(n320), .Z(n3166) );
  OAI21_X1 U2644 ( .B1(n4188), .B2(n4081), .A(n364), .ZN(n3911) );
  INV_X1 U2645 ( .A(n3911), .ZN(n3943) );
  MUX2_X1 U2646 ( .A(n4398), .B(n1033), .S(n321), .Z(n3912) );
  INV_X1 U2647 ( .A(n3912), .ZN(n3167) );
  MUX2_X1 U2648 ( .A(n4400), .B(n1074), .S(n321), .Z(n3913) );
  INV_X1 U2649 ( .A(n3913), .ZN(n3168) );
  MUX2_X1 U2650 ( .A(n4402), .B(n1110), .S(n321), .Z(n3914) );
  INV_X1 U2651 ( .A(n3914), .ZN(n3169) );
  MUX2_X1 U2652 ( .A(n4404), .B(n1146), .S(n321), .Z(n3915) );
  INV_X1 U2653 ( .A(n3915), .ZN(n3170) );
  MUX2_X1 U2654 ( .A(n4406), .B(n1182), .S(n321), .Z(n3916) );
  INV_X1 U2655 ( .A(n3916), .ZN(n3171) );
  MUX2_X1 U2656 ( .A(n4408), .B(n1218), .S(n321), .Z(n3917) );
  INV_X1 U2657 ( .A(n3917), .ZN(n3172) );
  MUX2_X1 U2658 ( .A(n4410), .B(n1254), .S(n321), .Z(n3918) );
  INV_X1 U2659 ( .A(n3918), .ZN(n3173) );
  MUX2_X1 U2660 ( .A(n4412), .B(n1290), .S(n321), .Z(n3919) );
  INV_X1 U2661 ( .A(n3919), .ZN(n3174) );
  MUX2_X1 U2662 ( .A(n4414), .B(n1326), .S(n321), .Z(n3920) );
  INV_X1 U2663 ( .A(n3920), .ZN(n3175) );
  MUX2_X1 U2664 ( .A(n4416), .B(n1362), .S(n321), .Z(n3921) );
  INV_X1 U2665 ( .A(n3921), .ZN(n3176) );
  MUX2_X1 U2666 ( .A(n4418), .B(n1398), .S(n321), .Z(n3922) );
  INV_X1 U2667 ( .A(n3922), .ZN(n3177) );
  MUX2_X1 U2668 ( .A(n4420), .B(n1434), .S(n321), .Z(n3923) );
  INV_X1 U2669 ( .A(n3923), .ZN(n3178) );
  MUX2_X1 U2670 ( .A(n4422), .B(n1470), .S(n322), .Z(n3924) );
  INV_X1 U2671 ( .A(n3924), .ZN(n3179) );
  MUX2_X1 U2672 ( .A(n4424), .B(n1506), .S(n322), .Z(n3925) );
  INV_X1 U2673 ( .A(n3925), .ZN(n3180) );
  MUX2_X1 U2674 ( .A(n4426), .B(n1542), .S(n322), .Z(n3926) );
  INV_X1 U2675 ( .A(n3926), .ZN(n3181) );
  MUX2_X1 U2676 ( .A(n4428), .B(n1578), .S(n322), .Z(n3927) );
  INV_X1 U2677 ( .A(n3927), .ZN(n3182) );
  MUX2_X1 U2678 ( .A(n4430), .B(n1614), .S(n322), .Z(n3928) );
  INV_X1 U2679 ( .A(n3928), .ZN(n3183) );
  MUX2_X1 U2680 ( .A(n4432), .B(n1650), .S(n322), .Z(n3929) );
  INV_X1 U2681 ( .A(n3929), .ZN(n3184) );
  MUX2_X1 U2682 ( .A(n4434), .B(n1686), .S(n322), .Z(n3930) );
  INV_X1 U2683 ( .A(n3930), .ZN(n3185) );
  MUX2_X1 U2684 ( .A(n4436), .B(n1722), .S(n322), .Z(n3931) );
  INV_X1 U2685 ( .A(n3931), .ZN(n3186) );
  MUX2_X1 U2686 ( .A(n4438), .B(n1758), .S(n322), .Z(n3932) );
  INV_X1 U2687 ( .A(n3932), .ZN(n3187) );
  MUX2_X1 U2688 ( .A(n4440), .B(n1794), .S(n322), .Z(n3933) );
  INV_X1 U2689 ( .A(n3933), .ZN(n3188) );
  MUX2_X1 U2690 ( .A(n4442), .B(n1830), .S(n322), .Z(n3934) );
  INV_X1 U2691 ( .A(n3934), .ZN(n3189) );
  MUX2_X1 U2692 ( .A(n4444), .B(n1866), .S(n322), .Z(n3935) );
  INV_X1 U2693 ( .A(n3935), .ZN(n3190) );
  MUX2_X1 U2694 ( .A(n4446), .B(n1902), .S(n323), .Z(n3936) );
  INV_X1 U2695 ( .A(n3936), .ZN(n3191) );
  MUX2_X1 U2696 ( .A(n4448), .B(n1938), .S(n323), .Z(n3937) );
  INV_X1 U2697 ( .A(n3937), .ZN(n3192) );
  MUX2_X1 U2698 ( .A(n4450), .B(n1974), .S(n323), .Z(n3938) );
  INV_X1 U2699 ( .A(n3938), .ZN(n3193) );
  MUX2_X1 U2700 ( .A(n4452), .B(n2010), .S(n323), .Z(n3939) );
  INV_X1 U2701 ( .A(n3939), .ZN(n3194) );
  MUX2_X1 U2702 ( .A(n4454), .B(n2046), .S(n323), .Z(n3940) );
  INV_X1 U2703 ( .A(n3940), .ZN(n3195) );
  MUX2_X1 U2704 ( .A(n4456), .B(n2082), .S(n323), .Z(n3941) );
  INV_X1 U2705 ( .A(n3941), .ZN(n3196) );
  MUX2_X1 U2706 ( .A(n4458), .B(n2118), .S(n323), .Z(n3942) );
  INV_X1 U2707 ( .A(n3942), .ZN(n3197) );
  MUX2_X1 U2708 ( .A(n4461), .B(n2155), .S(n323), .Z(n3944) );
  INV_X1 U2709 ( .A(n3944), .ZN(n3198) );
  OAI21_X1 U2710 ( .B1(n4223), .B2(n4081), .A(n364), .ZN(n3945) );
  INV_X1 U2711 ( .A(n3945), .ZN(n3977) );
  MUX2_X1 U2712 ( .A(n4398), .B(n1032), .S(n324), .Z(n3946) );
  INV_X1 U2713 ( .A(n3946), .ZN(n3199) );
  MUX2_X1 U2714 ( .A(n4400), .B(n1073), .S(n324), .Z(n3947) );
  INV_X1 U2715 ( .A(n3947), .ZN(n3200) );
  MUX2_X1 U2716 ( .A(n4402), .B(n1109), .S(n324), .Z(n3948) );
  INV_X1 U2717 ( .A(n3948), .ZN(n3201) );
  MUX2_X1 U2718 ( .A(n4404), .B(n1145), .S(n324), .Z(n3949) );
  INV_X1 U2719 ( .A(n3949), .ZN(n3202) );
  MUX2_X1 U2720 ( .A(n4406), .B(n1181), .S(n324), .Z(n3950) );
  INV_X1 U2721 ( .A(n3950), .ZN(n3203) );
  MUX2_X1 U2722 ( .A(n4408), .B(n1217), .S(n324), .Z(n3951) );
  INV_X1 U2723 ( .A(n3951), .ZN(n3204) );
  MUX2_X1 U2724 ( .A(n4410), .B(n1253), .S(n324), .Z(n3952) );
  INV_X1 U2725 ( .A(n3952), .ZN(n3205) );
  MUX2_X1 U2726 ( .A(n4412), .B(n1289), .S(n324), .Z(n3953) );
  INV_X1 U2727 ( .A(n3953), .ZN(n3206) );
  MUX2_X1 U2728 ( .A(n4414), .B(n1325), .S(n324), .Z(n3954) );
  INV_X1 U2729 ( .A(n3954), .ZN(n3207) );
  MUX2_X1 U2730 ( .A(n4416), .B(n1361), .S(n324), .Z(n3955) );
  INV_X1 U2731 ( .A(n3955), .ZN(n3208) );
  MUX2_X1 U2732 ( .A(n4418), .B(n1397), .S(n324), .Z(n3956) );
  INV_X1 U2733 ( .A(n3956), .ZN(n3209) );
  MUX2_X1 U2734 ( .A(n4420), .B(n1433), .S(n324), .Z(n3957) );
  INV_X1 U2735 ( .A(n3957), .ZN(n3210) );
  MUX2_X1 U2736 ( .A(n4422), .B(n1469), .S(n325), .Z(n3958) );
  INV_X1 U2737 ( .A(n3958), .ZN(n3211) );
  MUX2_X1 U2738 ( .A(n4424), .B(n1505), .S(n325), .Z(n3959) );
  INV_X1 U2739 ( .A(n3959), .ZN(n3212) );
  MUX2_X1 U2740 ( .A(n4426), .B(n1541), .S(n325), .Z(n3960) );
  INV_X1 U2741 ( .A(n3960), .ZN(n3213) );
  MUX2_X1 U2742 ( .A(n4428), .B(n1577), .S(n325), .Z(n3961) );
  INV_X1 U2743 ( .A(n3961), .ZN(n3214) );
  MUX2_X1 U2744 ( .A(n4430), .B(n1613), .S(n325), .Z(n3962) );
  INV_X1 U2745 ( .A(n3962), .ZN(n3215) );
  MUX2_X1 U2746 ( .A(n4432), .B(n1649), .S(n325), .Z(n3963) );
  INV_X1 U2747 ( .A(n3963), .ZN(n3216) );
  MUX2_X1 U2748 ( .A(n4434), .B(n1685), .S(n325), .Z(n3964) );
  INV_X1 U2749 ( .A(n3964), .ZN(n3217) );
  MUX2_X1 U2750 ( .A(n4436), .B(n1721), .S(n325), .Z(n3965) );
  INV_X1 U2751 ( .A(n3965), .ZN(n3218) );
  MUX2_X1 U2752 ( .A(n4438), .B(n1757), .S(n325), .Z(n3966) );
  INV_X1 U2753 ( .A(n3966), .ZN(n3219) );
  MUX2_X1 U2754 ( .A(n4440), .B(n1793), .S(n325), .Z(n3967) );
  INV_X1 U2755 ( .A(n3967), .ZN(n3220) );
  MUX2_X1 U2756 ( .A(n4442), .B(n1829), .S(n325), .Z(n3968) );
  INV_X1 U2757 ( .A(n3968), .ZN(n3221) );
  MUX2_X1 U2758 ( .A(n4444), .B(n1865), .S(n325), .Z(n3969) );
  INV_X1 U2759 ( .A(n3969), .ZN(n3222) );
  MUX2_X1 U2760 ( .A(n4446), .B(n1901), .S(n326), .Z(n3970) );
  INV_X1 U2761 ( .A(n3970), .ZN(n3223) );
  MUX2_X1 U2762 ( .A(n4448), .B(n1937), .S(n326), .Z(n3971) );
  INV_X1 U2763 ( .A(n3971), .ZN(n3224) );
  MUX2_X1 U2764 ( .A(n4450), .B(n1973), .S(n326), .Z(n3972) );
  INV_X1 U2765 ( .A(n3972), .ZN(n3225) );
  MUX2_X1 U2766 ( .A(n4452), .B(n2009), .S(n326), .Z(n3973) );
  INV_X1 U2767 ( .A(n3973), .ZN(n3226) );
  MUX2_X1 U2768 ( .A(n4454), .B(n2045), .S(n326), .Z(n3974) );
  INV_X1 U2769 ( .A(n3974), .ZN(n3227) );
  MUX2_X1 U2770 ( .A(n4456), .B(n2081), .S(n326), .Z(n3975) );
  INV_X1 U2771 ( .A(n3975), .ZN(n3228) );
  MUX2_X1 U2772 ( .A(n4458), .B(n2117), .S(n326), .Z(n3976) );
  INV_X1 U2773 ( .A(n3976), .ZN(n3229) );
  MUX2_X1 U2774 ( .A(n4461), .B(n2153), .S(n326), .Z(n3978) );
  INV_X1 U2775 ( .A(n3978), .ZN(n3230) );
  OAI21_X1 U2776 ( .B1(n4258), .B2(n4081), .A(n363), .ZN(n3979) );
  INV_X1 U2777 ( .A(n3979), .ZN(n4011) );
  MUX2_X1 U2778 ( .A(n4296), .B(n3980), .S(n327), .Z(n3231) );
  MUX2_X1 U2779 ( .A(n4298), .B(n3981), .S(n327), .Z(n3232) );
  MUX2_X1 U2780 ( .A(n4300), .B(n3982), .S(n327), .Z(n3233) );
  MUX2_X1 U2781 ( .A(n4302), .B(n3983), .S(n327), .Z(n3234) );
  MUX2_X1 U2782 ( .A(n4304), .B(n3984), .S(n327), .Z(n3235) );
  MUX2_X1 U2783 ( .A(n4306), .B(n3985), .S(n327), .Z(n3236) );
  MUX2_X1 U2784 ( .A(n4308), .B(n3986), .S(n327), .Z(n3237) );
  MUX2_X1 U2785 ( .A(n4310), .B(n3987), .S(n327), .Z(n3238) );
  MUX2_X1 U2786 ( .A(n4312), .B(n3988), .S(n327), .Z(n3239) );
  MUX2_X1 U2787 ( .A(n4314), .B(n3989), .S(n327), .Z(n3240) );
  MUX2_X1 U2788 ( .A(n4316), .B(n3990), .S(n327), .Z(n3241) );
  MUX2_X1 U2789 ( .A(n4318), .B(n3991), .S(n327), .Z(n3242) );
  MUX2_X1 U2790 ( .A(n4320), .B(n3992), .S(n328), .Z(n3243) );
  MUX2_X1 U2791 ( .A(n4322), .B(n3993), .S(n328), .Z(n3244) );
  MUX2_X1 U2792 ( .A(n4324), .B(n3994), .S(n328), .Z(n3245) );
  MUX2_X1 U2793 ( .A(n4326), .B(n3995), .S(n328), .Z(n3246) );
  MUX2_X1 U2794 ( .A(n4328), .B(n3996), .S(n328), .Z(n3247) );
  MUX2_X1 U2795 ( .A(n4330), .B(n3997), .S(n328), .Z(n3248) );
  MUX2_X1 U2796 ( .A(n4332), .B(n3998), .S(n328), .Z(n3249) );
  MUX2_X1 U2797 ( .A(n4334), .B(n3999), .S(n328), .Z(n3250) );
  MUX2_X1 U2798 ( .A(n4336), .B(n4000), .S(n328), .Z(n3251) );
  MUX2_X1 U2799 ( .A(n4338), .B(n4001), .S(n328), .Z(n3252) );
  MUX2_X1 U2800 ( .A(n4340), .B(n4002), .S(n328), .Z(n3253) );
  MUX2_X1 U2801 ( .A(n4342), .B(n4003), .S(n328), .Z(n3254) );
  MUX2_X1 U2802 ( .A(n4344), .B(n4004), .S(n329), .Z(n3255) );
  MUX2_X1 U2803 ( .A(n4346), .B(n4005), .S(n329), .Z(n3256) );
  MUX2_X1 U2804 ( .A(n4348), .B(n4006), .S(n329), .Z(n3257) );
  MUX2_X1 U2805 ( .A(n4350), .B(n4007), .S(n329), .Z(n3258) );
  MUX2_X1 U2806 ( .A(n4352), .B(n4008), .S(n329), .Z(n3259) );
  MUX2_X1 U2807 ( .A(n4354), .B(n4009), .S(n329), .Z(n3260) );
  MUX2_X1 U2808 ( .A(n4356), .B(n4010), .S(n329), .Z(n3261) );
  MUX2_X1 U2809 ( .A(n4359), .B(n4012), .S(n329), .Z(n3262) );
  OAI21_X1 U2810 ( .B1(n4293), .B2(n4081), .A(n363), .ZN(n4013) );
  INV_X1 U2811 ( .A(n4013), .ZN(n4045) );
  MUX2_X1 U2812 ( .A(n4296), .B(n4014), .S(n330), .Z(n3263) );
  MUX2_X1 U2813 ( .A(n4298), .B(n4015), .S(n330), .Z(n3264) );
  MUX2_X1 U2814 ( .A(n4300), .B(n4016), .S(n330), .Z(n3265) );
  MUX2_X1 U2815 ( .A(n4302), .B(n4017), .S(n330), .Z(n3266) );
  MUX2_X1 U2816 ( .A(n4304), .B(n4018), .S(n330), .Z(n3267) );
  MUX2_X1 U2817 ( .A(n4306), .B(n4019), .S(n330), .Z(n3268) );
  MUX2_X1 U2818 ( .A(n4308), .B(n4020), .S(n330), .Z(n3269) );
  MUX2_X1 U2819 ( .A(n4310), .B(n4021), .S(n330), .Z(n3270) );
  MUX2_X1 U2820 ( .A(n4312), .B(n4022), .S(n330), .Z(n3271) );
  MUX2_X1 U2821 ( .A(n4314), .B(n4023), .S(n330), .Z(n3272) );
  MUX2_X1 U2822 ( .A(n4316), .B(n4024), .S(n330), .Z(n3273) );
  MUX2_X1 U2823 ( .A(n4318), .B(n4025), .S(n330), .Z(n3274) );
  MUX2_X1 U2824 ( .A(n4320), .B(n4026), .S(n331), .Z(n3275) );
  MUX2_X1 U2825 ( .A(n4322), .B(n4027), .S(n331), .Z(n3276) );
  MUX2_X1 U2826 ( .A(n4324), .B(n4028), .S(n331), .Z(n3277) );
  MUX2_X1 U2827 ( .A(n4326), .B(n4029), .S(n331), .Z(n3278) );
  MUX2_X1 U2828 ( .A(n4328), .B(n4030), .S(n331), .Z(n3279) );
  MUX2_X1 U2829 ( .A(n4330), .B(n4031), .S(n331), .Z(n3280) );
  MUX2_X1 U2830 ( .A(n4332), .B(n4032), .S(n331), .Z(n3281) );
  MUX2_X1 U2831 ( .A(n4334), .B(n4033), .S(n331), .Z(n3282) );
  MUX2_X1 U2832 ( .A(n4336), .B(n4034), .S(n331), .Z(n3283) );
  MUX2_X1 U2833 ( .A(n4338), .B(n4035), .S(n331), .Z(n3284) );
  MUX2_X1 U2834 ( .A(n4340), .B(n4036), .S(n331), .Z(n3285) );
  MUX2_X1 U2835 ( .A(n4342), .B(n4037), .S(n331), .Z(n3286) );
  MUX2_X1 U2836 ( .A(n4344), .B(n4038), .S(n332), .Z(n3287) );
  MUX2_X1 U2837 ( .A(n4346), .B(n4039), .S(n332), .Z(n3288) );
  MUX2_X1 U2838 ( .A(n4348), .B(n4040), .S(n332), .Z(n3289) );
  MUX2_X1 U2839 ( .A(n4350), .B(n4041), .S(n332), .Z(n3290) );
  MUX2_X1 U2840 ( .A(n4352), .B(n4042), .S(n332), .Z(n3291) );
  MUX2_X1 U2841 ( .A(n4354), .B(n4043), .S(n332), .Z(n3292) );
  MUX2_X1 U2842 ( .A(n4356), .B(n4044), .S(n332), .Z(n3293) );
  MUX2_X1 U2843 ( .A(n4359), .B(n4046), .S(n332), .Z(n3294) );
  OAI21_X1 U2844 ( .B1(n4360), .B2(n4081), .A(n363), .ZN(n4047) );
  INV_X1 U2845 ( .A(n4047), .ZN(n4079) );
  MUX2_X1 U2846 ( .A(n4398), .B(n1038), .S(n333), .Z(n4048) );
  INV_X1 U2847 ( .A(n4048), .ZN(n3295) );
  MUX2_X1 U2848 ( .A(n4400), .B(n1077), .S(n333), .Z(n4049) );
  INV_X1 U2849 ( .A(n4049), .ZN(n3296) );
  MUX2_X1 U2850 ( .A(n4402), .B(n1113), .S(n333), .Z(n4050) );
  INV_X1 U2851 ( .A(n4050), .ZN(n3297) );
  MUX2_X1 U2852 ( .A(n4404), .B(n1149), .S(n333), .Z(n4051) );
  INV_X1 U2853 ( .A(n4051), .ZN(n3298) );
  MUX2_X1 U2854 ( .A(n4406), .B(n1185), .S(n333), .Z(n4052) );
  INV_X1 U2855 ( .A(n4052), .ZN(n3299) );
  MUX2_X1 U2856 ( .A(n4408), .B(n1221), .S(n333), .Z(n4053) );
  INV_X1 U2857 ( .A(n4053), .ZN(n3300) );
  MUX2_X1 U2858 ( .A(n4410), .B(n1257), .S(n333), .Z(n4054) );
  INV_X1 U2859 ( .A(n4054), .ZN(n3301) );
  MUX2_X1 U2860 ( .A(n4412), .B(n1293), .S(n333), .Z(n4055) );
  INV_X1 U2861 ( .A(n4055), .ZN(n3302) );
  MUX2_X1 U2862 ( .A(n4414), .B(n1329), .S(n333), .Z(n4056) );
  INV_X1 U2863 ( .A(n4056), .ZN(n3303) );
  MUX2_X1 U2864 ( .A(n4416), .B(n1365), .S(n333), .Z(n4057) );
  INV_X1 U2865 ( .A(n4057), .ZN(n3304) );
  MUX2_X1 U2866 ( .A(n4418), .B(n1401), .S(n333), .Z(n4058) );
  INV_X1 U2867 ( .A(n4058), .ZN(n3305) );
  MUX2_X1 U2868 ( .A(n4420), .B(n1437), .S(n333), .Z(n4059) );
  INV_X1 U2869 ( .A(n4059), .ZN(n3306) );
  MUX2_X1 U2870 ( .A(n4422), .B(n1473), .S(n334), .Z(n4060) );
  INV_X1 U2871 ( .A(n4060), .ZN(n3307) );
  MUX2_X1 U2872 ( .A(n4424), .B(n1509), .S(n334), .Z(n4061) );
  INV_X1 U2873 ( .A(n4061), .ZN(n3308) );
  MUX2_X1 U2874 ( .A(n4426), .B(n1545), .S(n334), .Z(n4062) );
  INV_X1 U2875 ( .A(n4062), .ZN(n3309) );
  MUX2_X1 U2876 ( .A(n4428), .B(n1581), .S(n334), .Z(n4063) );
  INV_X1 U2877 ( .A(n4063), .ZN(n3310) );
  MUX2_X1 U2878 ( .A(n4430), .B(n1617), .S(n334), .Z(n4064) );
  INV_X1 U2879 ( .A(n4064), .ZN(n3311) );
  MUX2_X1 U2880 ( .A(n4432), .B(n1653), .S(n334), .Z(n4065) );
  INV_X1 U2881 ( .A(n4065), .ZN(n3312) );
  MUX2_X1 U2882 ( .A(n4434), .B(n1689), .S(n334), .Z(n4066) );
  INV_X1 U2883 ( .A(n4066), .ZN(n3313) );
  MUX2_X1 U2884 ( .A(n4436), .B(n1725), .S(n334), .Z(n4067) );
  INV_X1 U2885 ( .A(n4067), .ZN(n3314) );
  MUX2_X1 U2886 ( .A(n4438), .B(n1761), .S(n334), .Z(n4068) );
  INV_X1 U2887 ( .A(n4068), .ZN(n3315) );
  MUX2_X1 U2888 ( .A(n4440), .B(n1797), .S(n334), .Z(n4069) );
  INV_X1 U2889 ( .A(n4069), .ZN(n3316) );
  MUX2_X1 U2890 ( .A(n4442), .B(n1833), .S(n334), .Z(n4070) );
  INV_X1 U2891 ( .A(n4070), .ZN(n3317) );
  MUX2_X1 U2892 ( .A(n4444), .B(n1869), .S(n334), .Z(n4071) );
  INV_X1 U2893 ( .A(n4071), .ZN(n3318) );
  MUX2_X1 U2894 ( .A(n4446), .B(n1905), .S(n335), .Z(n4072) );
  INV_X1 U2895 ( .A(n4072), .ZN(n3319) );
  MUX2_X1 U2896 ( .A(n4448), .B(n1941), .S(n335), .Z(n4073) );
  INV_X1 U2897 ( .A(n4073), .ZN(n3320) );
  MUX2_X1 U2898 ( .A(n4450), .B(n1977), .S(n335), .Z(n4074) );
  INV_X1 U2899 ( .A(n4074), .ZN(n3321) );
  MUX2_X1 U2900 ( .A(n4452), .B(n2013), .S(n335), .Z(n4075) );
  INV_X1 U2901 ( .A(n4075), .ZN(n3322) );
  MUX2_X1 U2902 ( .A(n4454), .B(n2049), .S(n335), .Z(n4076) );
  INV_X1 U2903 ( .A(n4076), .ZN(n3323) );
  MUX2_X1 U2904 ( .A(n4456), .B(n2085), .S(n335), .Z(n4077) );
  INV_X1 U2905 ( .A(n4077), .ZN(n3324) );
  MUX2_X1 U2906 ( .A(n4458), .B(n2121), .S(n335), .Z(n4078) );
  INV_X1 U2907 ( .A(n4078), .ZN(n3325) );
  MUX2_X1 U2908 ( .A(n4461), .B(n2160), .S(n335), .Z(n4080) );
  INV_X1 U2909 ( .A(n4080), .ZN(n3326) );
  OAI21_X1 U2910 ( .B1(n4395), .B2(n4081), .A(n363), .ZN(n4082) );
  INV_X1 U2911 ( .A(n4082), .ZN(n4114) );
  MUX2_X1 U2912 ( .A(n4398), .B(n1037), .S(n336), .Z(n4083) );
  INV_X1 U2913 ( .A(n4083), .ZN(n3327) );
  MUX2_X1 U2914 ( .A(n4400), .B(n1076), .S(n336), .Z(n4084) );
  INV_X1 U2915 ( .A(n4084), .ZN(n3328) );
  MUX2_X1 U2916 ( .A(n4402), .B(n1112), .S(n336), .Z(n4085) );
  INV_X1 U2917 ( .A(n4085), .ZN(n3329) );
  MUX2_X1 U2918 ( .A(n4404), .B(n1148), .S(n336), .Z(n4086) );
  INV_X1 U2919 ( .A(n4086), .ZN(n3330) );
  MUX2_X1 U2920 ( .A(n4406), .B(n1184), .S(n336), .Z(n4087) );
  INV_X1 U2921 ( .A(n4087), .ZN(n3331) );
  MUX2_X1 U2922 ( .A(n4408), .B(n1220), .S(n336), .Z(n4088) );
  INV_X1 U2923 ( .A(n4088), .ZN(n3332) );
  MUX2_X1 U2924 ( .A(n4410), .B(n1256), .S(n336), .Z(n4089) );
  INV_X1 U2925 ( .A(n4089), .ZN(n3333) );
  MUX2_X1 U2926 ( .A(n4412), .B(n1292), .S(n336), .Z(n4090) );
  INV_X1 U2927 ( .A(n4090), .ZN(n3334) );
  MUX2_X1 U2928 ( .A(n4414), .B(n1328), .S(n336), .Z(n4091) );
  INV_X1 U2929 ( .A(n4091), .ZN(n3335) );
  MUX2_X1 U2930 ( .A(n4416), .B(n1364), .S(n336), .Z(n4092) );
  INV_X1 U2931 ( .A(n4092), .ZN(n3336) );
  MUX2_X1 U2932 ( .A(n4418), .B(n1400), .S(n336), .Z(n4093) );
  INV_X1 U2933 ( .A(n4093), .ZN(n3337) );
  MUX2_X1 U2934 ( .A(n4420), .B(n1436), .S(n336), .Z(n4094) );
  INV_X1 U2935 ( .A(n4094), .ZN(n3338) );
  MUX2_X1 U2936 ( .A(n4422), .B(n1472), .S(n337), .Z(n4095) );
  INV_X1 U2937 ( .A(n4095), .ZN(n3339) );
  MUX2_X1 U2938 ( .A(n4424), .B(n1508), .S(n337), .Z(n4096) );
  INV_X1 U2939 ( .A(n4096), .ZN(n3340) );
  MUX2_X1 U2940 ( .A(n4426), .B(n1544), .S(n337), .Z(n4097) );
  INV_X1 U2941 ( .A(n4097), .ZN(n3341) );
  MUX2_X1 U2942 ( .A(n4428), .B(n1580), .S(n337), .Z(n4098) );
  INV_X1 U2943 ( .A(n4098), .ZN(n3342) );
  MUX2_X1 U2944 ( .A(n4430), .B(n1616), .S(n337), .Z(n4099) );
  INV_X1 U2945 ( .A(n4099), .ZN(n3343) );
  MUX2_X1 U2946 ( .A(n4432), .B(n1652), .S(n337), .Z(n4100) );
  INV_X1 U2947 ( .A(n4100), .ZN(n3344) );
  MUX2_X1 U2948 ( .A(n4434), .B(n1688), .S(n337), .Z(n4101) );
  INV_X1 U2949 ( .A(n4101), .ZN(n3345) );
  MUX2_X1 U2950 ( .A(n4436), .B(n1724), .S(n337), .Z(n4102) );
  INV_X1 U2951 ( .A(n4102), .ZN(n3346) );
  MUX2_X1 U2952 ( .A(n4438), .B(n1760), .S(n337), .Z(n4103) );
  INV_X1 U2953 ( .A(n4103), .ZN(n3347) );
  MUX2_X1 U2954 ( .A(n4440), .B(n1796), .S(n337), .Z(n4104) );
  INV_X1 U2955 ( .A(n4104), .ZN(n3348) );
  MUX2_X1 U2956 ( .A(n4442), .B(n1832), .S(n337), .Z(n4105) );
  INV_X1 U2957 ( .A(n4105), .ZN(n3349) );
  MUX2_X1 U2958 ( .A(n4444), .B(n1868), .S(n337), .Z(n4106) );
  INV_X1 U2959 ( .A(n4106), .ZN(n3350) );
  MUX2_X1 U2960 ( .A(n4446), .B(n1904), .S(n338), .Z(n4107) );
  INV_X1 U2961 ( .A(n4107), .ZN(n3351) );
  MUX2_X1 U2962 ( .A(n4448), .B(n1940), .S(n338), .Z(n4108) );
  INV_X1 U2963 ( .A(n4108), .ZN(n3352) );
  MUX2_X1 U2964 ( .A(n4450), .B(n1976), .S(n338), .Z(n4109) );
  INV_X1 U2965 ( .A(n4109), .ZN(n3353) );
  MUX2_X1 U2966 ( .A(n4452), .B(n2012), .S(n338), .Z(n4110) );
  INV_X1 U2967 ( .A(n4110), .ZN(n3354) );
  MUX2_X1 U2968 ( .A(n4454), .B(n2048), .S(n338), .Z(n4111) );
  INV_X1 U2969 ( .A(n4111), .ZN(n3355) );
  MUX2_X1 U2970 ( .A(n4456), .B(n2084), .S(n338), .Z(n4112) );
  INV_X1 U2971 ( .A(n4112), .ZN(n3356) );
  MUX2_X1 U2972 ( .A(n4458), .B(n2120), .S(n338), .Z(n4113) );
  INV_X1 U2973 ( .A(n4113), .ZN(n3357) );
  MUX2_X1 U2974 ( .A(n4461), .B(n2158), .S(n338), .Z(n4115) );
  INV_X1 U2975 ( .A(n4115), .ZN(n3358) );
  NAND3_X1 U2976 ( .A1(WR), .A2(n4117), .A3(n4116), .ZN(n4396) );
  OAI21_X1 U2977 ( .B1(n4396), .B2(n4118), .A(n363), .ZN(n4119) );
  INV_X1 U2978 ( .A(n4119), .ZN(n4151) );
  MUX2_X1 U2979 ( .A(n4296), .B(n4120), .S(n339), .Z(n3359) );
  MUX2_X1 U2980 ( .A(n4298), .B(n4121), .S(n339), .Z(n3360) );
  MUX2_X1 U2981 ( .A(n4300), .B(n4122), .S(n339), .Z(n3361) );
  MUX2_X1 U2982 ( .A(n4302), .B(n4123), .S(n339), .Z(n3362) );
  MUX2_X1 U2983 ( .A(n4304), .B(n4124), .S(n339), .Z(n3363) );
  MUX2_X1 U2984 ( .A(n4306), .B(n4125), .S(n339), .Z(n3364) );
  MUX2_X1 U2985 ( .A(n4308), .B(n4126), .S(n339), .Z(n3365) );
  MUX2_X1 U2986 ( .A(n4310), .B(n4127), .S(n339), .Z(n3366) );
  MUX2_X1 U2987 ( .A(n4312), .B(n4128), .S(n339), .Z(n3367) );
  MUX2_X1 U2988 ( .A(n4314), .B(n4129), .S(n339), .Z(n3368) );
  MUX2_X1 U2989 ( .A(n4316), .B(n4130), .S(n339), .Z(n3369) );
  MUX2_X1 U2990 ( .A(n4318), .B(n4131), .S(n339), .Z(n3370) );
  MUX2_X1 U2991 ( .A(n4320), .B(n4132), .S(n340), .Z(n3371) );
  MUX2_X1 U2992 ( .A(n4322), .B(n4133), .S(n340), .Z(n3372) );
  MUX2_X1 U2993 ( .A(n4324), .B(n4134), .S(n340), .Z(n3373) );
  MUX2_X1 U2994 ( .A(n4326), .B(n4135), .S(n340), .Z(n3374) );
  MUX2_X1 U2995 ( .A(n4328), .B(n4136), .S(n340), .Z(n3375) );
  MUX2_X1 U2996 ( .A(n4330), .B(n4137), .S(n340), .Z(n3376) );
  MUX2_X1 U2997 ( .A(n4332), .B(n4138), .S(n340), .Z(n3377) );
  MUX2_X1 U2998 ( .A(n4334), .B(n4139), .S(n340), .Z(n3378) );
  MUX2_X1 U2999 ( .A(n4336), .B(n4140), .S(n340), .Z(n3379) );
  MUX2_X1 U3000 ( .A(n4338), .B(n4141), .S(n340), .Z(n3380) );
  MUX2_X1 U3001 ( .A(n4340), .B(n4142), .S(n340), .Z(n3381) );
  MUX2_X1 U3002 ( .A(n4342), .B(n4143), .S(n340), .Z(n3382) );
  MUX2_X1 U3003 ( .A(n4344), .B(n4144), .S(n341), .Z(n3383) );
  MUX2_X1 U3004 ( .A(n4346), .B(n4145), .S(n341), .Z(n3384) );
  MUX2_X1 U3005 ( .A(n4348), .B(n4146), .S(n341), .Z(n3385) );
  MUX2_X1 U3006 ( .A(n4350), .B(n4147), .S(n341), .Z(n3386) );
  MUX2_X1 U3007 ( .A(n4352), .B(n4148), .S(n341), .Z(n3387) );
  MUX2_X1 U3008 ( .A(n4354), .B(n4149), .S(n341), .Z(n3388) );
  MUX2_X1 U3009 ( .A(n4356), .B(n4150), .S(n341), .Z(n3389) );
  MUX2_X1 U3010 ( .A(n4359), .B(n4152), .S(n341), .Z(n3390) );
  OAI21_X1 U3011 ( .B1(n4396), .B2(n4153), .A(n363), .ZN(n4154) );
  INV_X1 U3012 ( .A(n4154), .ZN(n4186) );
  MUX2_X1 U3013 ( .A(n4296), .B(n4155), .S(n342), .Z(n3391) );
  MUX2_X1 U3014 ( .A(n4298), .B(n4156), .S(n342), .Z(n3392) );
  MUX2_X1 U3015 ( .A(n4300), .B(n4157), .S(n342), .Z(n3393) );
  MUX2_X1 U3016 ( .A(n4302), .B(n4158), .S(n342), .Z(n3394) );
  MUX2_X1 U3017 ( .A(n4304), .B(n4159), .S(n342), .Z(n3395) );
  MUX2_X1 U3018 ( .A(n4306), .B(n4160), .S(n342), .Z(n3396) );
  MUX2_X1 U3019 ( .A(n4308), .B(n4161), .S(n342), .Z(n3397) );
  MUX2_X1 U3020 ( .A(n4310), .B(n4162), .S(n342), .Z(n3398) );
  MUX2_X1 U3021 ( .A(n4312), .B(n4163), .S(n342), .Z(n3399) );
  MUX2_X1 U3022 ( .A(n4314), .B(n4164), .S(n342), .Z(n3400) );
  MUX2_X1 U3023 ( .A(n4316), .B(n4165), .S(n342), .Z(n3401) );
  MUX2_X1 U3024 ( .A(n4318), .B(n4166), .S(n342), .Z(n3402) );
  MUX2_X1 U3025 ( .A(n4320), .B(n4167), .S(n343), .Z(n3403) );
  MUX2_X1 U3026 ( .A(n4322), .B(n4168), .S(n343), .Z(n3404) );
  MUX2_X1 U3027 ( .A(n4324), .B(n4169), .S(n343), .Z(n3405) );
  MUX2_X1 U3028 ( .A(n4326), .B(n4170), .S(n343), .Z(n3406) );
  MUX2_X1 U3029 ( .A(n4328), .B(n4171), .S(n343), .Z(n3407) );
  MUX2_X1 U3030 ( .A(n4330), .B(n4172), .S(n343), .Z(n3408) );
  MUX2_X1 U3031 ( .A(n4332), .B(n4173), .S(n343), .Z(n3409) );
  MUX2_X1 U3032 ( .A(n4334), .B(n4174), .S(n343), .Z(n3410) );
  MUX2_X1 U3033 ( .A(n4336), .B(n4175), .S(n343), .Z(n3411) );
  MUX2_X1 U3034 ( .A(n4338), .B(n4176), .S(n343), .Z(n3412) );
  MUX2_X1 U3035 ( .A(n4340), .B(n4177), .S(n343), .Z(n3413) );
  MUX2_X1 U3036 ( .A(n4342), .B(n4178), .S(n343), .Z(n3414) );
  MUX2_X1 U3037 ( .A(n4344), .B(n4179), .S(n344), .Z(n3415) );
  MUX2_X1 U3038 ( .A(n4346), .B(n4180), .S(n344), .Z(n3416) );
  MUX2_X1 U3039 ( .A(n4348), .B(n4181), .S(n344), .Z(n3417) );
  MUX2_X1 U3040 ( .A(n4350), .B(n4182), .S(n344), .Z(n3418) );
  MUX2_X1 U3041 ( .A(n4352), .B(n4183), .S(n344), .Z(n3419) );
  MUX2_X1 U3042 ( .A(n4354), .B(n4184), .S(n344), .Z(n3420) );
  MUX2_X1 U3043 ( .A(n4356), .B(n4185), .S(n344), .Z(n3421) );
  MUX2_X1 U3044 ( .A(n4359), .B(n4187), .S(n344), .Z(n3422) );
  OAI21_X1 U3045 ( .B1(n4396), .B2(n4188), .A(n363), .ZN(n4189) );
  INV_X1 U3046 ( .A(n4189), .ZN(n4221) );
  MUX2_X1 U3047 ( .A(n4398), .B(n1042), .S(n345), .Z(n4190) );
  INV_X1 U3048 ( .A(n4190), .ZN(n3423) );
  MUX2_X1 U3049 ( .A(n4400), .B(n1080), .S(n345), .Z(n4191) );
  INV_X1 U3050 ( .A(n4191), .ZN(n3424) );
  MUX2_X1 U3051 ( .A(n4402), .B(n1116), .S(n345), .Z(n4192) );
  INV_X1 U3052 ( .A(n4192), .ZN(n3425) );
  MUX2_X1 U3053 ( .A(n4404), .B(n1152), .S(n345), .Z(n4193) );
  INV_X1 U3054 ( .A(n4193), .ZN(n3426) );
  MUX2_X1 U3055 ( .A(n4406), .B(n1188), .S(n345), .Z(n4194) );
  INV_X1 U3056 ( .A(n4194), .ZN(n3427) );
  MUX2_X1 U3057 ( .A(n4408), .B(n1224), .S(n345), .Z(n4195) );
  INV_X1 U3058 ( .A(n4195), .ZN(n3428) );
  MUX2_X1 U3059 ( .A(n4410), .B(n1260), .S(n345), .Z(n4196) );
  INV_X1 U3060 ( .A(n4196), .ZN(n3429) );
  MUX2_X1 U3061 ( .A(n4412), .B(n1296), .S(n345), .Z(n4197) );
  INV_X1 U3062 ( .A(n4197), .ZN(n3430) );
  MUX2_X1 U3063 ( .A(n4414), .B(n1332), .S(n345), .Z(n4198) );
  INV_X1 U3064 ( .A(n4198), .ZN(n3431) );
  MUX2_X1 U3065 ( .A(n4416), .B(n1368), .S(n345), .Z(n4199) );
  INV_X1 U3066 ( .A(n4199), .ZN(n3432) );
  MUX2_X1 U3067 ( .A(n4418), .B(n1404), .S(n345), .Z(n4200) );
  INV_X1 U3068 ( .A(n4200), .ZN(n3433) );
  MUX2_X1 U3069 ( .A(n4420), .B(n1440), .S(n345), .Z(n4201) );
  INV_X1 U3070 ( .A(n4201), .ZN(n3434) );
  MUX2_X1 U3071 ( .A(n4422), .B(n1476), .S(n346), .Z(n4202) );
  INV_X1 U3072 ( .A(n4202), .ZN(n3435) );
  MUX2_X1 U3073 ( .A(n4424), .B(n1512), .S(n346), .Z(n4203) );
  INV_X1 U3074 ( .A(n4203), .ZN(n3436) );
  MUX2_X1 U3075 ( .A(n4426), .B(n1548), .S(n346), .Z(n4204) );
  INV_X1 U3076 ( .A(n4204), .ZN(n3437) );
  MUX2_X1 U3077 ( .A(n4428), .B(n1584), .S(n346), .Z(n4205) );
  INV_X1 U3078 ( .A(n4205), .ZN(n3438) );
  MUX2_X1 U3079 ( .A(n4430), .B(n1620), .S(n346), .Z(n4206) );
  INV_X1 U3080 ( .A(n4206), .ZN(n3439) );
  MUX2_X1 U3081 ( .A(n4432), .B(n1656), .S(n346), .Z(n4207) );
  INV_X1 U3082 ( .A(n4207), .ZN(n3440) );
  MUX2_X1 U3083 ( .A(n4434), .B(n1692), .S(n346), .Z(n4208) );
  INV_X1 U3084 ( .A(n4208), .ZN(n3441) );
  MUX2_X1 U3085 ( .A(n4436), .B(n1728), .S(n346), .Z(n4209) );
  INV_X1 U3086 ( .A(n4209), .ZN(n3442) );
  MUX2_X1 U3087 ( .A(n4438), .B(n1764), .S(n346), .Z(n4210) );
  INV_X1 U3088 ( .A(n4210), .ZN(n3443) );
  MUX2_X1 U3089 ( .A(n4440), .B(n1800), .S(n346), .Z(n4211) );
  INV_X1 U3090 ( .A(n4211), .ZN(n3444) );
  MUX2_X1 U3091 ( .A(n4442), .B(n1836), .S(n346), .Z(n4212) );
  INV_X1 U3092 ( .A(n4212), .ZN(n3445) );
  MUX2_X1 U3093 ( .A(n4444), .B(n1872), .S(n346), .Z(n4213) );
  INV_X1 U3094 ( .A(n4213), .ZN(n3446) );
  MUX2_X1 U3095 ( .A(n4446), .B(n1908), .S(n347), .Z(n4214) );
  INV_X1 U3096 ( .A(n4214), .ZN(n3447) );
  MUX2_X1 U3097 ( .A(n4448), .B(n1944), .S(n347), .Z(n4215) );
  INV_X1 U3098 ( .A(n4215), .ZN(n3448) );
  MUX2_X1 U3099 ( .A(n4450), .B(n1980), .S(n347), .Z(n4216) );
  INV_X1 U3100 ( .A(n4216), .ZN(n3449) );
  MUX2_X1 U3101 ( .A(n4452), .B(n2016), .S(n347), .Z(n4217) );
  INV_X1 U3102 ( .A(n4217), .ZN(n3450) );
  MUX2_X1 U3103 ( .A(n4454), .B(n2052), .S(n347), .Z(n4218) );
  INV_X1 U3104 ( .A(n4218), .ZN(n3451) );
  MUX2_X1 U3105 ( .A(n4456), .B(n2088), .S(n347), .Z(n4219) );
  INV_X1 U3106 ( .A(n4219), .ZN(n3452) );
  MUX2_X1 U3107 ( .A(n4458), .B(n2124), .S(n347), .Z(n4220) );
  INV_X1 U3108 ( .A(n4220), .ZN(n3453) );
  MUX2_X1 U3109 ( .A(n4461), .B(n2165), .S(n347), .Z(n4222) );
  INV_X1 U3110 ( .A(n4222), .ZN(n3454) );
  OAI21_X1 U3111 ( .B1(n4396), .B2(n4223), .A(n363), .ZN(n4224) );
  INV_X1 U3112 ( .A(n4224), .ZN(n4256) );
  MUX2_X1 U3113 ( .A(n4398), .B(n1041), .S(n348), .Z(n4225) );
  INV_X1 U3114 ( .A(n4225), .ZN(n3455) );
  MUX2_X1 U3115 ( .A(n4400), .B(n1079), .S(n348), .Z(n4226) );
  INV_X1 U3116 ( .A(n4226), .ZN(n3456) );
  MUX2_X1 U3117 ( .A(n4402), .B(n1115), .S(n348), .Z(n4227) );
  INV_X1 U3118 ( .A(n4227), .ZN(n3457) );
  MUX2_X1 U3119 ( .A(n4404), .B(n1151), .S(n348), .Z(n4228) );
  INV_X1 U3120 ( .A(n4228), .ZN(n3458) );
  MUX2_X1 U3121 ( .A(n4406), .B(n1187), .S(n348), .Z(n4229) );
  INV_X1 U3122 ( .A(n4229), .ZN(n3459) );
  MUX2_X1 U3123 ( .A(n4408), .B(n1223), .S(n348), .Z(n4230) );
  INV_X1 U3124 ( .A(n4230), .ZN(n3460) );
  MUX2_X1 U3125 ( .A(n4410), .B(n1259), .S(n348), .Z(n4231) );
  INV_X1 U3126 ( .A(n4231), .ZN(n3461) );
  MUX2_X1 U3127 ( .A(n4412), .B(n1295), .S(n348), .Z(n4232) );
  INV_X1 U3128 ( .A(n4232), .ZN(n3462) );
  MUX2_X1 U3129 ( .A(n4414), .B(n1331), .S(n348), .Z(n4233) );
  INV_X1 U3130 ( .A(n4233), .ZN(n3463) );
  MUX2_X1 U3131 ( .A(n4416), .B(n1367), .S(n348), .Z(n4234) );
  INV_X1 U3132 ( .A(n4234), .ZN(n3464) );
  MUX2_X1 U3133 ( .A(n4418), .B(n1403), .S(n348), .Z(n4235) );
  INV_X1 U3134 ( .A(n4235), .ZN(n3465) );
  MUX2_X1 U3135 ( .A(n4420), .B(n1439), .S(n348), .Z(n4236) );
  INV_X1 U3136 ( .A(n4236), .ZN(n3466) );
  MUX2_X1 U3137 ( .A(n4422), .B(n1475), .S(n349), .Z(n4237) );
  INV_X1 U3138 ( .A(n4237), .ZN(n3467) );
  MUX2_X1 U3139 ( .A(n4424), .B(n1511), .S(n349), .Z(n4238) );
  INV_X1 U3140 ( .A(n4238), .ZN(n3468) );
  MUX2_X1 U3141 ( .A(n4426), .B(n1547), .S(n349), .Z(n4239) );
  INV_X1 U3142 ( .A(n4239), .ZN(n3469) );
  MUX2_X1 U3143 ( .A(n4428), .B(n1583), .S(n349), .Z(n4240) );
  INV_X1 U3144 ( .A(n4240), .ZN(n3470) );
  MUX2_X1 U3145 ( .A(n4430), .B(n1619), .S(n349), .Z(n4241) );
  INV_X1 U3146 ( .A(n4241), .ZN(n3471) );
  MUX2_X1 U3147 ( .A(n4432), .B(n1655), .S(n349), .Z(n4242) );
  INV_X1 U3148 ( .A(n4242), .ZN(n3472) );
  MUX2_X1 U3149 ( .A(n4434), .B(n1691), .S(n349), .Z(n4243) );
  INV_X1 U3150 ( .A(n4243), .ZN(n3473) );
  MUX2_X1 U3151 ( .A(n4436), .B(n1727), .S(n349), .Z(n4244) );
  INV_X1 U3152 ( .A(n4244), .ZN(n3474) );
  MUX2_X1 U3153 ( .A(n4438), .B(n1763), .S(n349), .Z(n4245) );
  INV_X1 U3154 ( .A(n4245), .ZN(n3475) );
  MUX2_X1 U3155 ( .A(n4440), .B(n1799), .S(n349), .Z(n4246) );
  INV_X1 U3156 ( .A(n4246), .ZN(n3476) );
  MUX2_X1 U3157 ( .A(n4442), .B(n1835), .S(n349), .Z(n4247) );
  INV_X1 U3158 ( .A(n4247), .ZN(n3477) );
  MUX2_X1 U3159 ( .A(n4444), .B(n1871), .S(n349), .Z(n4248) );
  INV_X1 U3160 ( .A(n4248), .ZN(n3478) );
  MUX2_X1 U3161 ( .A(n4446), .B(n1907), .S(n350), .Z(n4249) );
  INV_X1 U3162 ( .A(n4249), .ZN(n3479) );
  MUX2_X1 U3163 ( .A(n4448), .B(n1943), .S(n350), .Z(n4250) );
  INV_X1 U3164 ( .A(n4250), .ZN(n3480) );
  MUX2_X1 U3165 ( .A(n4450), .B(n1979), .S(n350), .Z(n4251) );
  INV_X1 U3166 ( .A(n4251), .ZN(n3481) );
  MUX2_X1 U3167 ( .A(n4452), .B(n2015), .S(n350), .Z(n4252) );
  INV_X1 U3168 ( .A(n4252), .ZN(n3482) );
  MUX2_X1 U3169 ( .A(n4454), .B(n2051), .S(n350), .Z(n4253) );
  INV_X1 U3170 ( .A(n4253), .ZN(n3483) );
  MUX2_X1 U3171 ( .A(n4456), .B(n2087), .S(n350), .Z(n4254) );
  INV_X1 U3172 ( .A(n4254), .ZN(n3484) );
  MUX2_X1 U3173 ( .A(n4458), .B(n2123), .S(n350), .Z(n4255) );
  INV_X1 U3174 ( .A(n4255), .ZN(n3485) );
  MUX2_X1 U3175 ( .A(n4461), .B(n2163), .S(n350), .Z(n4257) );
  INV_X1 U3176 ( .A(n4257), .ZN(n3486) );
  OAI21_X1 U3177 ( .B1(n4396), .B2(n4258), .A(n363), .ZN(n4259) );
  INV_X1 U3178 ( .A(n4259), .ZN(n4291) );
  MUX2_X1 U3179 ( .A(n4296), .B(n4260), .S(n351), .Z(n3487) );
  MUX2_X1 U3180 ( .A(n4298), .B(n4261), .S(n351), .Z(n3488) );
  MUX2_X1 U3181 ( .A(n4300), .B(n4262), .S(n351), .Z(n3489) );
  MUX2_X1 U3182 ( .A(n4302), .B(n4263), .S(n351), .Z(n3490) );
  MUX2_X1 U3183 ( .A(n4304), .B(n4264), .S(n351), .Z(n3491) );
  MUX2_X1 U3184 ( .A(n4306), .B(n4265), .S(n351), .Z(n3492) );
  MUX2_X1 U3185 ( .A(n4308), .B(n4266), .S(n351), .Z(n3493) );
  MUX2_X1 U3186 ( .A(n4310), .B(n4267), .S(n351), .Z(n3494) );
  MUX2_X1 U3187 ( .A(n4312), .B(n4268), .S(n351), .Z(n3495) );
  MUX2_X1 U3188 ( .A(n4314), .B(n4269), .S(n351), .Z(n3496) );
  MUX2_X1 U3189 ( .A(n4316), .B(n4270), .S(n351), .Z(n3497) );
  MUX2_X1 U3190 ( .A(n4318), .B(n4271), .S(n351), .Z(n3498) );
  MUX2_X1 U3191 ( .A(n4320), .B(n4272), .S(n352), .Z(n3499) );
  MUX2_X1 U3192 ( .A(n4322), .B(n4273), .S(n352), .Z(n3500) );
  MUX2_X1 U3193 ( .A(n4324), .B(n4274), .S(n352), .Z(n3501) );
  MUX2_X1 U3194 ( .A(n4326), .B(n4275), .S(n352), .Z(n3502) );
  MUX2_X1 U3195 ( .A(n4328), .B(n4276), .S(n352), .Z(n3503) );
  MUX2_X1 U3196 ( .A(n4330), .B(n4277), .S(n352), .Z(n3504) );
  MUX2_X1 U3197 ( .A(n4332), .B(n4278), .S(n352), .Z(n3505) );
  MUX2_X1 U3198 ( .A(n4334), .B(n4279), .S(n352), .Z(n3506) );
  MUX2_X1 U3199 ( .A(n4336), .B(n4280), .S(n352), .Z(n3507) );
  MUX2_X1 U3200 ( .A(n4338), .B(n4281), .S(n352), .Z(n3508) );
  MUX2_X1 U3201 ( .A(n4340), .B(n4282), .S(n352), .Z(n3509) );
  MUX2_X1 U3202 ( .A(n4342), .B(n4283), .S(n352), .Z(n3510) );
  MUX2_X1 U3203 ( .A(n4344), .B(n4284), .S(n353), .Z(n3511) );
  MUX2_X1 U3204 ( .A(n4346), .B(n4285), .S(n353), .Z(n3512) );
  MUX2_X1 U3205 ( .A(n4348), .B(n4286), .S(n353), .Z(n3513) );
  MUX2_X1 U3206 ( .A(n4350), .B(n4287), .S(n353), .Z(n3514) );
  MUX2_X1 U3207 ( .A(n4352), .B(n4288), .S(n353), .Z(n3515) );
  MUX2_X1 U3208 ( .A(n4354), .B(n4289), .S(n353), .Z(n3516) );
  MUX2_X1 U3209 ( .A(n4356), .B(n4290), .S(n353), .Z(n3517) );
  MUX2_X1 U3210 ( .A(n4359), .B(n4292), .S(n353), .Z(n3518) );
  OAI21_X1 U3211 ( .B1(n4396), .B2(n4293), .A(n363), .ZN(n4294) );
  INV_X1 U3212 ( .A(n4294), .ZN(n4357) );
  MUX2_X1 U3213 ( .A(n4296), .B(n4295), .S(n354), .Z(n3519) );
  MUX2_X1 U3214 ( .A(n4298), .B(n4297), .S(n354), .Z(n3520) );
  MUX2_X1 U3215 ( .A(n4300), .B(n4299), .S(n354), .Z(n3521) );
  MUX2_X1 U3216 ( .A(n4302), .B(n4301), .S(n354), .Z(n3522) );
  MUX2_X1 U3217 ( .A(n4304), .B(n4303), .S(n354), .Z(n3523) );
  MUX2_X1 U3218 ( .A(n4306), .B(n4305), .S(n354), .Z(n3524) );
  MUX2_X1 U3219 ( .A(n4308), .B(n4307), .S(n354), .Z(n3525) );
  MUX2_X1 U3220 ( .A(n4310), .B(n4309), .S(n354), .Z(n3526) );
  MUX2_X1 U3221 ( .A(n4312), .B(n4311), .S(n354), .Z(n3527) );
  MUX2_X1 U3222 ( .A(n4314), .B(n4313), .S(n354), .Z(n3528) );
  MUX2_X1 U3223 ( .A(n4316), .B(n4315), .S(n354), .Z(n3529) );
  MUX2_X1 U3224 ( .A(n4318), .B(n4317), .S(n354), .Z(n3530) );
  MUX2_X1 U3225 ( .A(n4320), .B(n4319), .S(n355), .Z(n3531) );
  MUX2_X1 U3226 ( .A(n4322), .B(n4321), .S(n355), .Z(n3532) );
  MUX2_X1 U3227 ( .A(n4324), .B(n4323), .S(n355), .Z(n3533) );
  MUX2_X1 U3228 ( .A(n4326), .B(n4325), .S(n355), .Z(n3534) );
  MUX2_X1 U3229 ( .A(n4328), .B(n4327), .S(n355), .Z(n3535) );
  MUX2_X1 U3230 ( .A(n4330), .B(n4329), .S(n355), .Z(n3536) );
  MUX2_X1 U3231 ( .A(n4332), .B(n4331), .S(n355), .Z(n3537) );
  MUX2_X1 U3232 ( .A(n4334), .B(n4333), .S(n355), .Z(n3538) );
  MUX2_X1 U3233 ( .A(n4336), .B(n4335), .S(n355), .Z(n3539) );
  MUX2_X1 U3234 ( .A(n4338), .B(n4337), .S(n355), .Z(n3540) );
  MUX2_X1 U3235 ( .A(n4340), .B(n4339), .S(n355), .Z(n3541) );
  MUX2_X1 U3236 ( .A(n4342), .B(n4341), .S(n355), .Z(n3542) );
  MUX2_X1 U3237 ( .A(n4344), .B(n4343), .S(n356), .Z(n3543) );
  MUX2_X1 U3238 ( .A(n4346), .B(n4345), .S(n356), .Z(n3544) );
  MUX2_X1 U3239 ( .A(n4348), .B(n4347), .S(n356), .Z(n3545) );
  MUX2_X1 U3240 ( .A(n4350), .B(n4349), .S(n356), .Z(n3546) );
  MUX2_X1 U3241 ( .A(n4352), .B(n4351), .S(n356), .Z(n3547) );
  MUX2_X1 U3242 ( .A(n4354), .B(n4353), .S(n356), .Z(n3548) );
  MUX2_X1 U3243 ( .A(n4356), .B(n4355), .S(n356), .Z(n3549) );
  MUX2_X1 U3244 ( .A(n4359), .B(n4358), .S(n356), .Z(n3550) );
  OAI21_X1 U3245 ( .B1(n4396), .B2(n4360), .A(n363), .ZN(n4361) );
  INV_X1 U3246 ( .A(n4361), .ZN(n4393) );
  MUX2_X1 U3247 ( .A(n4398), .B(n1045), .S(n357), .Z(n4362) );
  INV_X1 U3248 ( .A(n4362), .ZN(n3551) );
  MUX2_X1 U3249 ( .A(n4400), .B(n1083), .S(n357), .Z(n4363) );
  INV_X1 U3250 ( .A(n4363), .ZN(n3552) );
  MUX2_X1 U3251 ( .A(n4402), .B(n1119), .S(n357), .Z(n4364) );
  INV_X1 U3252 ( .A(n4364), .ZN(n3553) );
  MUX2_X1 U3253 ( .A(n4404), .B(n1155), .S(n357), .Z(n4365) );
  INV_X1 U3254 ( .A(n4365), .ZN(n3554) );
  MUX2_X1 U3255 ( .A(n4406), .B(n1191), .S(n357), .Z(n4366) );
  INV_X1 U3256 ( .A(n4366), .ZN(n3555) );
  MUX2_X1 U3257 ( .A(n4408), .B(n1227), .S(n357), .Z(n4367) );
  INV_X1 U3258 ( .A(n4367), .ZN(n3556) );
  MUX2_X1 U3259 ( .A(n4410), .B(n1263), .S(n357), .Z(n4368) );
  INV_X1 U3260 ( .A(n4368), .ZN(n3557) );
  MUX2_X1 U3261 ( .A(n4412), .B(n1299), .S(n357), .Z(n4369) );
  INV_X1 U3262 ( .A(n4369), .ZN(n3558) );
  MUX2_X1 U3263 ( .A(n4414), .B(n1335), .S(n357), .Z(n4370) );
  INV_X1 U3264 ( .A(n4370), .ZN(n3559) );
  MUX2_X1 U3265 ( .A(n4416), .B(n1371), .S(n357), .Z(n4371) );
  INV_X1 U3266 ( .A(n4371), .ZN(n3560) );
  MUX2_X1 U3267 ( .A(n4418), .B(n1407), .S(n357), .Z(n4372) );
  INV_X1 U3268 ( .A(n4372), .ZN(n3561) );
  MUX2_X1 U3269 ( .A(n4420), .B(n1443), .S(n357), .Z(n4373) );
  INV_X1 U3270 ( .A(n4373), .ZN(n3562) );
  MUX2_X1 U3271 ( .A(n4422), .B(n1479), .S(n358), .Z(n4374) );
  INV_X1 U3272 ( .A(n4374), .ZN(n3563) );
  MUX2_X1 U3273 ( .A(n4424), .B(n1515), .S(n358), .Z(n4375) );
  INV_X1 U3274 ( .A(n4375), .ZN(n3564) );
  MUX2_X1 U3275 ( .A(n4426), .B(n1551), .S(n358), .Z(n4376) );
  INV_X1 U3276 ( .A(n4376), .ZN(n3565) );
  MUX2_X1 U3277 ( .A(n4428), .B(n1587), .S(n358), .Z(n4377) );
  INV_X1 U3278 ( .A(n4377), .ZN(n3566) );
  MUX2_X1 U3279 ( .A(n4430), .B(n1623), .S(n358), .Z(n4378) );
  INV_X1 U3280 ( .A(n4378), .ZN(n3567) );
  MUX2_X1 U3281 ( .A(n4432), .B(n1659), .S(n358), .Z(n4379) );
  INV_X1 U3282 ( .A(n4379), .ZN(n3568) );
  MUX2_X1 U3283 ( .A(n4434), .B(n1695), .S(n358), .Z(n4380) );
  INV_X1 U3284 ( .A(n4380), .ZN(n3569) );
  MUX2_X1 U3285 ( .A(n4436), .B(n1731), .S(n358), .Z(n4381) );
  INV_X1 U3286 ( .A(n4381), .ZN(n3570) );
  MUX2_X1 U3287 ( .A(n4438), .B(n1767), .S(n358), .Z(n4382) );
  INV_X1 U3288 ( .A(n4382), .ZN(n3571) );
  MUX2_X1 U3289 ( .A(n4440), .B(n1803), .S(n358), .Z(n4383) );
  INV_X1 U3290 ( .A(n4383), .ZN(n3572) );
  MUX2_X1 U3291 ( .A(n4442), .B(n1839), .S(n358), .Z(n4384) );
  INV_X1 U3292 ( .A(n4384), .ZN(n3573) );
  MUX2_X1 U3293 ( .A(n4444), .B(n1875), .S(n358), .Z(n4385) );
  INV_X1 U3294 ( .A(n4385), .ZN(n3574) );
  MUX2_X1 U3295 ( .A(n4446), .B(n1911), .S(n359), .Z(n4386) );
  INV_X1 U3296 ( .A(n4386), .ZN(n3575) );
  MUX2_X1 U3297 ( .A(n4448), .B(n1947), .S(n359), .Z(n4387) );
  INV_X1 U3298 ( .A(n4387), .ZN(n3576) );
  MUX2_X1 U3299 ( .A(n4450), .B(n1983), .S(n359), .Z(n4388) );
  INV_X1 U3300 ( .A(n4388), .ZN(n3577) );
  MUX2_X1 U3301 ( .A(n4452), .B(n2019), .S(n359), .Z(n4389) );
  INV_X1 U3302 ( .A(n4389), .ZN(n3578) );
  MUX2_X1 U3303 ( .A(n4454), .B(n2055), .S(n359), .Z(n4390) );
  INV_X1 U3304 ( .A(n4390), .ZN(n3579) );
  MUX2_X1 U3305 ( .A(n4456), .B(n2091), .S(n359), .Z(n4391) );
  INV_X1 U3306 ( .A(n4391), .ZN(n3580) );
  MUX2_X1 U3307 ( .A(n4458), .B(n2127), .S(n359), .Z(n4392) );
  INV_X1 U3308 ( .A(n4392), .ZN(n3581) );
  MUX2_X1 U3309 ( .A(n4461), .B(n2170), .S(n359), .Z(n4394) );
  INV_X1 U3310 ( .A(n4394), .ZN(n3582) );
  OAI21_X1 U3311 ( .B1(n4396), .B2(n4395), .A(n364), .ZN(n4397) );
  INV_X1 U3312 ( .A(n4397), .ZN(n4460) );
  MUX2_X1 U3313 ( .A(n4398), .B(n1044), .S(n360), .Z(n4399) );
  INV_X1 U3314 ( .A(n4399), .ZN(n3583) );
  MUX2_X1 U3315 ( .A(n4400), .B(n1082), .S(n360), .Z(n4401) );
  INV_X1 U3316 ( .A(n4401), .ZN(n3584) );
  MUX2_X1 U3317 ( .A(n4402), .B(n1118), .S(n360), .Z(n4403) );
  INV_X1 U3318 ( .A(n4403), .ZN(n3585) );
  MUX2_X1 U3319 ( .A(n4404), .B(n1154), .S(n360), .Z(n4405) );
  INV_X1 U3320 ( .A(n4405), .ZN(n3586) );
  MUX2_X1 U3321 ( .A(n4406), .B(n1190), .S(n360), .Z(n4407) );
  INV_X1 U3322 ( .A(n4407), .ZN(n3587) );
  MUX2_X1 U3323 ( .A(n4408), .B(n1226), .S(n360), .Z(n4409) );
  INV_X1 U3324 ( .A(n4409), .ZN(n3588) );
  MUX2_X1 U3325 ( .A(n4410), .B(n1262), .S(n360), .Z(n4411) );
  INV_X1 U3326 ( .A(n4411), .ZN(n3589) );
  MUX2_X1 U3327 ( .A(n4412), .B(n1298), .S(n360), .Z(n4413) );
  INV_X1 U3328 ( .A(n4413), .ZN(n3590) );
  MUX2_X1 U3329 ( .A(n4414), .B(n1334), .S(n360), .Z(n4415) );
  INV_X1 U3330 ( .A(n4415), .ZN(n3591) );
  MUX2_X1 U3331 ( .A(n4416), .B(n1370), .S(n360), .Z(n4417) );
  INV_X1 U3332 ( .A(n4417), .ZN(n3592) );
  MUX2_X1 U3333 ( .A(n4418), .B(n1406), .S(n360), .Z(n4419) );
  INV_X1 U3334 ( .A(n4419), .ZN(n3593) );
  MUX2_X1 U3335 ( .A(n4420), .B(n1442), .S(n360), .Z(n4421) );
  INV_X1 U3336 ( .A(n4421), .ZN(n3594) );
  MUX2_X1 U3337 ( .A(n4422), .B(n1478), .S(n361), .Z(n4423) );
  INV_X1 U3338 ( .A(n4423), .ZN(n3595) );
  MUX2_X1 U3339 ( .A(n4424), .B(n1514), .S(n361), .Z(n4425) );
  INV_X1 U3340 ( .A(n4425), .ZN(n3596) );
  MUX2_X1 U3341 ( .A(n4426), .B(n1550), .S(n361), .Z(n4427) );
  INV_X1 U3342 ( .A(n4427), .ZN(n3597) );
  MUX2_X1 U3343 ( .A(n4428), .B(n1586), .S(n361), .Z(n4429) );
  INV_X1 U3344 ( .A(n4429), .ZN(n3598) );
  MUX2_X1 U3345 ( .A(n4430), .B(n1622), .S(n361), .Z(n4431) );
  INV_X1 U3346 ( .A(n4431), .ZN(n3599) );
  MUX2_X1 U3347 ( .A(n4432), .B(n1658), .S(n361), .Z(n4433) );
  INV_X1 U3348 ( .A(n4433), .ZN(n3600) );
  MUX2_X1 U3349 ( .A(n4434), .B(n1694), .S(n361), .Z(n4435) );
  INV_X1 U3350 ( .A(n4435), .ZN(n3601) );
  MUX2_X1 U3351 ( .A(n4436), .B(n1730), .S(n361), .Z(n4437) );
  INV_X1 U3352 ( .A(n4437), .ZN(n3602) );
  MUX2_X1 U3353 ( .A(n4438), .B(n1766), .S(n361), .Z(n4439) );
  INV_X1 U3354 ( .A(n4439), .ZN(n3603) );
  MUX2_X1 U3355 ( .A(n4440), .B(n1802), .S(n361), .Z(n4441) );
  INV_X1 U3356 ( .A(n4441), .ZN(n3604) );
  MUX2_X1 U3357 ( .A(n4442), .B(n1838), .S(n361), .Z(n4443) );
  INV_X1 U3358 ( .A(n4443), .ZN(n3605) );
  MUX2_X1 U3359 ( .A(n4444), .B(n1874), .S(n361), .Z(n4445) );
  INV_X1 U3360 ( .A(n4445), .ZN(n3606) );
  MUX2_X1 U3361 ( .A(n4446), .B(n1910), .S(n362), .Z(n4447) );
  INV_X1 U3362 ( .A(n4447), .ZN(n3607) );
  MUX2_X1 U3363 ( .A(n4448), .B(n1946), .S(n362), .Z(n4449) );
  INV_X1 U3364 ( .A(n4449), .ZN(n3608) );
  MUX2_X1 U3365 ( .A(n4450), .B(n1982), .S(n362), .Z(n4451) );
  INV_X1 U3366 ( .A(n4451), .ZN(n3609) );
  MUX2_X1 U3367 ( .A(n4452), .B(n2018), .S(n362), .Z(n4453) );
  INV_X1 U3368 ( .A(n4453), .ZN(n3610) );
  MUX2_X1 U3369 ( .A(n4454), .B(n2054), .S(n362), .Z(n4455) );
  INV_X1 U3370 ( .A(n4455), .ZN(n3611) );
  MUX2_X1 U3371 ( .A(n4456), .B(n2090), .S(n362), .Z(n4457) );
  INV_X1 U3372 ( .A(n4457), .ZN(n3612) );
  MUX2_X1 U3373 ( .A(n4458), .B(n2126), .S(n362), .Z(n4459) );
  INV_X1 U3374 ( .A(n4459), .ZN(n3613) );
  MUX2_X1 U3375 ( .A(n4461), .B(n2168), .S(n362), .Z(n4462) );
  INV_X1 U3376 ( .A(n4462), .ZN(n3614) );
  DFF_X1 \OUT1_reg[31]  ( .D(n2590), .CK(CLK), .Q(OUT1[31]), .QN(n2204) );
  DFF_X1 \OUT1_reg[30]  ( .D(n2589), .CK(CLK), .Q(OUT1[30]), .QN(n2152) );
  DFF_X1 \OUT1_reg[29]  ( .D(n2588), .CK(CLK), .Q(OUT1[29]), .QN(n2116) );
  DFF_X1 \OUT1_reg[28]  ( .D(n2587), .CK(CLK), .Q(OUT1[28]), .QN(n2080) );
  DFF_X1 \OUT1_reg[27]  ( .D(n2586), .CK(CLK), .Q(OUT1[27]), .QN(n2044) );
  DFF_X1 \OUT1_reg[26]  ( .D(n2585), .CK(CLK), .Q(OUT1[26]), .QN(n2008) );
  DFF_X1 \OUT1_reg[25]  ( .D(n2584), .CK(CLK), .Q(OUT1[25]), .QN(n1972) );
  DFF_X1 \OUT1_reg[24]  ( .D(n2583), .CK(CLK), .Q(OUT1[24]), .QN(n1936) );
  DFF_X1 \OUT2_reg[31]  ( .D(n2558), .CK(CLK), .Q(OUT2[31]), .QN(n1030) );
  DFF_X1 \OUT2_reg[30]  ( .D(n2557), .CK(CLK), .Q(OUT2[30]), .QN(n994) );
  DFF_X1 \OUT2_reg[29]  ( .D(n2556), .CK(CLK), .Q(OUT2[29]), .QN(n974) );
  DFF_X1 \OUT2_reg[28]  ( .D(n2555), .CK(CLK), .Q(OUT2[28]), .QN(n954) );
  DFF_X1 \OUT2_reg[27]  ( .D(n2554), .CK(CLK), .Q(OUT2[27]), .QN(n934) );
  DFF_X1 \OUT2_reg[26]  ( .D(n2553), .CK(CLK), .Q(OUT2[26]), .QN(n914) );
  DFF_X1 \OUT2_reg[25]  ( .D(n2552), .CK(CLK), .Q(OUT2[25]), .QN(n894) );
  DFF_X1 \OUT2_reg[24]  ( .D(n2551), .CK(CLK), .Q(OUT2[24]), .QN(n874) );
  DFF_X1 \OUT1_reg[10]  ( .D(n2569), .CK(CLK), .Q(OUT1[10]), .QN(n1432) );
  DFF_X1 \OUT1_reg[9]  ( .D(n2568), .CK(CLK), .Q(OUT1[9]), .QN(n1396) );
  DFF_X1 \OUT1_reg[8]  ( .D(n2567), .CK(CLK), .Q(OUT1[8]), .QN(n1360) );
  DFF_X1 \OUT1_reg[7]  ( .D(n2566), .CK(CLK), .Q(OUT1[7]), .QN(n1324) );
  DFF_X1 \OUT1_reg[6]  ( .D(n2565), .CK(CLK), .Q(OUT1[6]), .QN(n1288) );
  DFF_X1 \OUT1_reg[5]  ( .D(n2564), .CK(CLK), .Q(OUT1[5]), .QN(n1252) );
  DFF_X1 \OUT1_reg[4]  ( .D(n2563), .CK(CLK), .Q(OUT1[4]), .QN(n1216) );
  DFF_X1 \OUT1_reg[3]  ( .D(n2562), .CK(CLK), .Q(OUT1[3]), .QN(n1180) );
  DFF_X1 \OUT1_reg[2]  ( .D(n2561), .CK(CLK), .Q(OUT1[2]), .QN(n1144) );
  DFF_X1 \OUT1_reg[1]  ( .D(n2560), .CK(CLK), .Q(OUT1[1]), .QN(n1108) );
  DFF_X1 \OUT1_reg[0]  ( .D(n2559), .CK(CLK), .Q(OUT1[0]), .QN(n1072) );
  DFF_X1 \OUT1_reg[23]  ( .D(n2582), .CK(CLK), .Q(OUT1[23]), .QN(n1900) );
  DFF_X1 \OUT1_reg[22]  ( .D(n2581), .CK(CLK), .Q(OUT1[22]), .QN(n1864) );
  DFF_X1 \OUT1_reg[21]  ( .D(n2580), .CK(CLK), .Q(OUT1[21]), .QN(n1828) );
  DFF_X1 \OUT1_reg[20]  ( .D(n2579), .CK(CLK), .Q(OUT1[20]), .QN(n1792) );
  DFF_X1 \OUT1_reg[19]  ( .D(n2578), .CK(CLK), .Q(OUT1[19]), .QN(n1756) );
  DFF_X1 \OUT1_reg[18]  ( .D(n2577), .CK(CLK), .Q(OUT1[18]), .QN(n1720) );
  DFF_X1 \OUT1_reg[17]  ( .D(n2576), .CK(CLK), .Q(OUT1[17]), .QN(n1684) );
  DFF_X1 \OUT1_reg[16]  ( .D(n2575), .CK(CLK), .Q(OUT1[16]), .QN(n1648) );
  DFF_X1 \OUT1_reg[15]  ( .D(n2574), .CK(CLK), .Q(OUT1[15]), .QN(n1612) );
  DFF_X1 \OUT1_reg[14]  ( .D(n2573), .CK(CLK), .Q(OUT1[14]), .QN(n1576) );
endmodule


module EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26 ( NOT_EXT_IMM, SIGNED_IMM, IS_JUMP, 
        EXT_IMM );
  input [25:0] NOT_EXT_IMM;
  output [31:0] EXT_IMM;
  input SIGNED_IMM, IS_JUMP;
  wire   \EXT_IMM[31] , \NOT_EXT_IMM[15] , \NOT_EXT_IMM[14] ,
         \NOT_EXT_IMM[13] , \NOT_EXT_IMM[12] , \NOT_EXT_IMM[11] ,
         \NOT_EXT_IMM[10] , \NOT_EXT_IMM[9] , \NOT_EXT_IMM[8] ,
         \NOT_EXT_IMM[7] , \NOT_EXT_IMM[6] , \NOT_EXT_IMM[5] ,
         \NOT_EXT_IMM[4] , \NOT_EXT_IMM[3] , \NOT_EXT_IMM[2] ,
         \NOT_EXT_IMM[1] , \NOT_EXT_IMM[0] , n2, n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23;
  assign EXT_IMM[26] = \EXT_IMM[31] ;
  assign EXT_IMM[27] = \EXT_IMM[31] ;
  assign EXT_IMM[28] = \EXT_IMM[31] ;
  assign EXT_IMM[29] = \EXT_IMM[31] ;
  assign EXT_IMM[30] = \EXT_IMM[31] ;
  assign EXT_IMM[31] = \EXT_IMM[31] ;
  assign EXT_IMM[15] = \NOT_EXT_IMM[15] ;
  assign \NOT_EXT_IMM[15]  = NOT_EXT_IMM[15];
  assign EXT_IMM[14] = \NOT_EXT_IMM[14] ;
  assign \NOT_EXT_IMM[14]  = NOT_EXT_IMM[14];
  assign EXT_IMM[13] = \NOT_EXT_IMM[13] ;
  assign \NOT_EXT_IMM[13]  = NOT_EXT_IMM[13];
  assign EXT_IMM[12] = \NOT_EXT_IMM[12] ;
  assign \NOT_EXT_IMM[12]  = NOT_EXT_IMM[12];
  assign EXT_IMM[11] = \NOT_EXT_IMM[11] ;
  assign \NOT_EXT_IMM[11]  = NOT_EXT_IMM[11];
  assign EXT_IMM[10] = \NOT_EXT_IMM[10] ;
  assign \NOT_EXT_IMM[10]  = NOT_EXT_IMM[10];
  assign EXT_IMM[9] = \NOT_EXT_IMM[9] ;
  assign \NOT_EXT_IMM[9]  = NOT_EXT_IMM[9];
  assign EXT_IMM[8] = \NOT_EXT_IMM[8] ;
  assign \NOT_EXT_IMM[8]  = NOT_EXT_IMM[8];
  assign EXT_IMM[7] = \NOT_EXT_IMM[7] ;
  assign \NOT_EXT_IMM[7]  = NOT_EXT_IMM[7];
  assign EXT_IMM[6] = \NOT_EXT_IMM[6] ;
  assign \NOT_EXT_IMM[6]  = NOT_EXT_IMM[6];
  assign EXT_IMM[5] = \NOT_EXT_IMM[5] ;
  assign \NOT_EXT_IMM[5]  = NOT_EXT_IMM[5];
  assign EXT_IMM[4] = \NOT_EXT_IMM[4] ;
  assign \NOT_EXT_IMM[4]  = NOT_EXT_IMM[4];
  assign EXT_IMM[3] = \NOT_EXT_IMM[3] ;
  assign \NOT_EXT_IMM[3]  = NOT_EXT_IMM[3];
  assign EXT_IMM[2] = \NOT_EXT_IMM[2] ;
  assign \NOT_EXT_IMM[2]  = NOT_EXT_IMM[2];
  assign EXT_IMM[1] = \NOT_EXT_IMM[1] ;
  assign \NOT_EXT_IMM[1]  = NOT_EXT_IMM[1];
  assign EXT_IMM[0] = \NOT_EXT_IMM[0] ;
  assign \NOT_EXT_IMM[0]  = NOT_EXT_IMM[0];

  OR2_X1 U2 ( .A1(n6), .A2(n18), .ZN(EXT_IMM[20]) );
  AND2_X1 U3 ( .A1(\NOT_EXT_IMM[15] ), .A2(SIGNED_IMM), .ZN(n2) );
  CLKBUF_X1 U4 ( .A(IS_JUMP), .Z(n3) );
  OR2_X1 U5 ( .A1(n7), .A2(n5), .ZN(EXT_IMM[18]) );
  AND3_X1 U6 ( .A1(\NOT_EXT_IMM[15] ), .A2(SIGNED_IMM), .A3(n22), .ZN(n5) );
  AND2_X1 U7 ( .A1(n9), .A2(NOT_EXT_IMM[20]), .ZN(n6) );
  AND2_X1 U8 ( .A1(n8), .A2(n2), .ZN(n10) );
  AND2_X1 U9 ( .A1(NOT_EXT_IMM[18]), .A2(n9), .ZN(n7) );
  INV_X1 U10 ( .A(IS_JUMP), .ZN(n8) );
  INV_X2 U11 ( .A(n8), .ZN(n9) );
  NAND2_X1 U12 ( .A1(n13), .A2(n12), .ZN(EXT_IMM[17]) );
  NAND2_X1 U13 ( .A1(NOT_EXT_IMM[17]), .A2(n3), .ZN(n12) );
  INV_X1 U14 ( .A(IS_JUMP), .ZN(n22) );
  NAND3_X1 U15 ( .A1(\NOT_EXT_IMM[15] ), .A2(n22), .A3(SIGNED_IMM), .ZN(n20)
         );
  INV_X1 U16 ( .A(n20), .ZN(n18) );
  AOI21_X1 U17 ( .B1(NOT_EXT_IMM[16]), .B2(n9), .A(n10), .ZN(n11) );
  INV_X1 U18 ( .A(n11), .ZN(EXT_IMM[16]) );
  NAND3_X1 U19 ( .A1(SIGNED_IMM), .A2(\NOT_EXT_IMM[15] ), .A3(n22), .ZN(n13)
         );
  AOI21_X1 U20 ( .B1(NOT_EXT_IMM[19]), .B2(n9), .A(n18), .ZN(n14) );
  INV_X1 U21 ( .A(n14), .ZN(EXT_IMM[19]) );
  AOI21_X1 U22 ( .B1(NOT_EXT_IMM[21]), .B2(n9), .A(n5), .ZN(n15) );
  INV_X1 U23 ( .A(n15), .ZN(EXT_IMM[21]) );
  AOI21_X1 U24 ( .B1(NOT_EXT_IMM[22]), .B2(n9), .A(n10), .ZN(n16) );
  INV_X1 U25 ( .A(n16), .ZN(EXT_IMM[22]) );
  AOI21_X1 U26 ( .B1(n9), .B2(NOT_EXT_IMM[23]), .A(n10), .ZN(n17) );
  INV_X1 U27 ( .A(n17), .ZN(EXT_IMM[23]) );
  AOI21_X1 U28 ( .B1(NOT_EXT_IMM[24]), .B2(n9), .A(n10), .ZN(n19) );
  INV_X1 U29 ( .A(n19), .ZN(EXT_IMM[24]) );
  INV_X1 U30 ( .A(NOT_EXT_IMM[25]), .ZN(n21) );
  OAI21_X1 U31 ( .B1(n22), .B2(n21), .A(n20), .ZN(EXT_IMM[25]) );
  OAI221_X1 U32 ( .B1(n8), .B2(NOT_EXT_IMM[25]), .C1(\NOT_EXT_IMM[15] ), .C2(
        n3), .A(SIGNED_IMM), .ZN(n23) );
  INV_X1 U33 ( .A(n23), .ZN(\EXT_IMM[31] ) );
endmodule


module NAND3_0 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_127 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_126 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_125 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_124 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_123 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_122 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_121 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_120 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_119 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_118 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_117 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_116 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_115 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_114 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_113 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_112 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_111 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_110 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_109 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_108 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_107 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_106 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_105 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_104 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_103 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_102 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_101 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_100 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_99 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_98 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_97 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_96 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_95 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_94 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_93 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_92 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_91 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_90 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_89 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_88 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_87 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_86 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_85 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_84 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_83 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_82 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_81 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_80 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_79 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_78 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_77 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_76 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_75 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_74 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_73 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_72 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_71 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_70 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_69 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_68 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_67 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_66 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_65 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_64 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_63 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_62 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_61 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_60 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_59 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_58 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_57 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_56 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_55 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_54 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_53 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_52 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_51 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_50 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_49 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_48 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_47 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_46 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_45 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_44 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_43 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_42 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_41 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_40 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_39 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_38 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_37 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_36 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_35 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_34 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_33 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_32 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_31 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_30 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_29 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_28 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_27 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_26 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_25 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_24 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_23 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_22 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_21 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_20 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_19 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_18 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_17 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_16 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_15 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_14 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_13 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_12 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_11 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_10 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_9 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_8 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_7 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_6 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_5 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_4 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_3 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_2 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND3_1 ( A, B, C, Y );
  input A, B, C;
  output Y;


  NAND3_X1 U1 ( .A1(B), .A2(A), .A3(C), .ZN(Y) );
endmodule


module NAND4_0 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_31 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_30 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_29 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_28 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_27 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_26 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_25 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_24 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_23 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_22 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_21 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_20 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_19 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_18 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_17 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_16 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_15 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_14 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_13 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_12 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_11 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_10 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_9 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_8 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_7 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_6 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_5 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_4 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_3 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_2 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module NAND4_1 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;


  NAND4_X1 U1 ( .A1(B), .A2(A), .A3(D), .A4(C), .ZN(Y) );
endmodule


module BARREL_SHIFTER_N32 ( CONF, DATA1, DATA2, OUTPUT );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUTPUT;
  input CONF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516;

  BUF_X1 U2 ( .A(n26), .Z(n16) );
  MUX2_X2 U3 ( .A(n443), .B(n418), .S(n138), .Z(n431) );
  CLKBUF_X3 U4 ( .A(n501), .Z(n37) );
  NAND3_X1 U5 ( .A1(n342), .A2(n112), .A3(n111), .ZN(n1) );
  CLKBUF_X1 U6 ( .A(DATA2[3]), .Z(n8) );
  INV_X1 U7 ( .A(n25), .ZN(n2) );
  MUX2_X1 U8 ( .A(n166), .B(n167), .S(n147), .Z(n174) );
  INV_X2 U9 ( .A(DATA2[2]), .ZN(n147) );
  NAND3_X1 U10 ( .A1(n61), .A2(n62), .A3(n190), .ZN(n3) );
  BUF_X2 U11 ( .A(n90), .Z(n115) );
  INV_X1 U12 ( .A(n313), .ZN(n4) );
  INV_X1 U13 ( .A(n355), .ZN(n5) );
  OR2_X1 U14 ( .A1(n69), .A2(n334), .ZN(n6) );
  OR2_X1 U15 ( .A1(n37), .A2(n414), .ZN(n7) );
  NAND3_X1 U16 ( .A1(n6), .A2(n7), .A3(n333), .ZN(n379) );
  CLKBUF_X1 U17 ( .A(DATA2[3]), .Z(n101) );
  AND3_X1 U18 ( .A1(n118), .A2(n332), .A3(n98), .ZN(n78) );
  OR3_X1 U19 ( .A1(n414), .A2(n8), .A3(n437), .ZN(n9) );
  OR2_X1 U20 ( .A1(n438), .A2(n8), .ZN(n10) );
  AOI221_X1 U21 ( .B1(n163), .B2(DATA1[16]), .C1(n162), .C2(DATA1[24]), .A(
        n148), .ZN(n152) );
  AND2_X1 U22 ( .A1(n103), .A2(n35), .ZN(n11) );
  NAND3_X1 U23 ( .A1(n43), .A2(n44), .A3(n391), .ZN(n12) );
  MUX2_X1 U24 ( .A(n249), .B(n259), .S(n133), .Z(n250) );
  INV_X1 U25 ( .A(n132), .ZN(n128) );
  NAND3_X1 U26 ( .A1(n67), .A2(n68), .A3(n185), .ZN(n13) );
  MUX2_X1 U27 ( .A(n18), .B(n19), .S(n147), .Z(n295) );
  INV_X1 U28 ( .A(n146), .ZN(n143) );
  NAND3_X1 U29 ( .A1(n65), .A2(n66), .A3(n199), .ZN(n14) );
  MUX2_X1 U30 ( .A(n233), .B(n216), .S(n140), .Z(n228) );
  INV_X2 U31 ( .A(n140), .ZN(n134) );
  OR2_X1 U32 ( .A1(n37), .A2(n343), .ZN(n15) );
  MUX2_X1 U33 ( .A(n296), .B(n278), .S(n135), .Z(n288) );
  NAND3_X1 U34 ( .A1(n15), .A2(n60), .A3(n266), .ZN(n17) );
  NAND3_X1 U35 ( .A1(n88), .A2(n89), .A3(n256), .ZN(n18) );
  NAND3_X1 U36 ( .A1(n294), .A2(n106), .A3(n105), .ZN(n19) );
  MUX2_X1 U37 ( .A(n336), .B(n346), .S(n132), .Z(n337) );
  MUX2_X1 U38 ( .A(n4), .B(n314), .S(n135), .Z(n20) );
  MUX2_X1 U39 ( .A(n434), .B(n1), .S(DATA2[2]), .Z(n384) );
  INV_X1 U40 ( .A(n282), .ZN(n21) );
  INV_X1 U41 ( .A(n313), .ZN(n22) );
  BUF_X2 U42 ( .A(n26), .Z(n23) );
  CLKBUF_X1 U43 ( .A(DATA1[7]), .Z(n24) );
  BUF_X2 U44 ( .A(n26), .Z(n113) );
  AND3_X2 U45 ( .A1(n332), .A2(n99), .A3(n125), .ZN(n26) );
  BUF_X2 U46 ( .A(n73), .Z(n25) );
  AND3_X1 U47 ( .A1(n332), .A2(n99), .A3(n125), .ZN(n90) );
  BUF_X1 U48 ( .A(n501), .Z(n108) );
  AND3_X1 U49 ( .A1(n332), .A2(n103), .A3(n118), .ZN(n27) );
  MUX2_X1 U50 ( .A(n22), .B(n356), .S(n140), .Z(n32) );
  MUX2_X1 U51 ( .A(n482), .B(n509), .S(n140), .Z(n494) );
  OR2_X1 U52 ( .A1(n83), .A2(n452), .ZN(n28) );
  OR2_X1 U53 ( .A1(n91), .A2(n451), .ZN(n29) );
  NAND3_X1 U54 ( .A1(n28), .A2(n29), .A3(n450), .ZN(n506) );
  MUX2_X1 U55 ( .A(n395), .B(n5), .S(n137), .Z(n30) );
  NAND3_X1 U56 ( .A1(n47), .A2(n48), .A3(n312), .ZN(n31) );
  MUX2_X1 U57 ( .A(n104), .B(n458), .S(n147), .Z(n406) );
  MUX2_X1 U58 ( .A(n430), .B(n407), .S(n134), .Z(n419) );
  NAND3_X1 U59 ( .A1(n383), .A2(n50), .A3(n49), .ZN(n33) );
  AOI221_X4 U60 ( .B1(n24), .B2(n41), .C1(DATA1[15]), .C2(n504), .A(n503), 
        .ZN(n508) );
  CLKBUF_X3 U61 ( .A(n116), .Z(n123) );
  OAI221_X1 U62 ( .B1(n83), .B2(n452), .C1(n91), .C2(n451), .A(n450), .ZN(n34)
         );
  NAND2_X1 U63 ( .A1(n103), .A2(n35), .ZN(n160) );
  AND2_X1 U64 ( .A1(DATA2[3]), .A2(n116), .ZN(n35) );
  CLKBUF_X1 U65 ( .A(CONF), .Z(n116) );
  MUX2_X1 U66 ( .A(n443), .B(n467), .S(n140), .Z(n455) );
  NAND2_X1 U67 ( .A1(n93), .A2(n100), .ZN(n36) );
  NAND2_X1 U68 ( .A1(n93), .A2(n100), .ZN(n246) );
  MUX2_X1 U69 ( .A(n431), .B(n444), .S(n133), .Z(n432) );
  INV_X1 U70 ( .A(n133), .ZN(n131) );
  MUX2_X1 U71 ( .A(n79), .B(n291), .S(n145), .Z(n286) );
  MUX2_X1 U72 ( .A(n305), .B(n325), .S(n140), .Z(n315) );
  INV_X1 U73 ( .A(n139), .ZN(n136) );
  INV_X2 U74 ( .A(DATA2[1]), .ZN(n140) );
  MUX2_X1 U75 ( .A(n418), .B(n395), .S(n137), .Z(n408) );
  MUX2_X1 U76 ( .A(n38), .B(n330), .S(n136), .Z(n321) );
  NOR2_X1 U77 ( .A1(n39), .A2(n40), .ZN(n38) );
  AND2_X1 U78 ( .A1(n328), .A2(n142), .ZN(n39) );
  AND2_X1 U79 ( .A1(n291), .A2(n92), .ZN(n40) );
  MUX2_X1 U80 ( .A(n14), .B(n291), .S(n147), .Z(n247) );
  INV_X2 U81 ( .A(n139), .ZN(n135) );
  INV_X2 U82 ( .A(n133), .ZN(n130) );
  INV_X1 U83 ( .A(n478), .ZN(n41) );
  INV_X1 U84 ( .A(n139), .ZN(n138) );
  CLKBUF_X3 U85 ( .A(n116), .Z(n122) );
  OAI221_X1 U86 ( .B1(n25), .B2(n393), .C1(n487), .C2(n36), .A(n235), .ZN(n42)
         );
  MUX2_X1 U87 ( .A(n318), .B(n42), .S(DATA2[2]), .Z(n277) );
  AOI22_X1 U88 ( .A1(n26), .A2(DATA1[31]), .B1(n27), .B2(DATA1[23]), .ZN(n403)
         );
  OR2_X1 U89 ( .A1(n91), .A2(n393), .ZN(n43) );
  OR2_X1 U90 ( .A1(n37), .A2(n392), .ZN(n44) );
  NAND3_X1 U91 ( .A1(n43), .A2(n44), .A3(n391), .ZN(n447) );
  NAND3_X1 U92 ( .A1(n51), .A2(n52), .A3(n374), .ZN(n45) );
  NAND3_X1 U93 ( .A1(n342), .A2(n112), .A3(n111), .ZN(n46) );
  INV_X1 U94 ( .A(n26), .ZN(n159) );
  MUX2_X1 U95 ( .A(n430), .B(n454), .S(n139), .Z(n444) );
  OR2_X1 U96 ( .A1(n108), .A2(n393), .ZN(n47) );
  OR2_X1 U97 ( .A1(n110), .A2(n392), .ZN(n48) );
  NAND3_X1 U98 ( .A1(n47), .A2(n48), .A3(n312), .ZN(n360) );
  OR2_X1 U99 ( .A1(n69), .A2(n477), .ZN(n49) );
  OR2_X1 U100 ( .A1(n37), .A2(n476), .ZN(n50) );
  NAND3_X1 U101 ( .A1(n49), .A2(n50), .A3(n383), .ZN(n434) );
  OR2_X1 U102 ( .A1(n91), .A2(n463), .ZN(n51) );
  OR2_X1 U103 ( .A1(n37), .A2(n462), .ZN(n52) );
  NAND3_X1 U104 ( .A1(n51), .A2(n52), .A3(n374), .ZN(n422) );
  OR2_X1 U105 ( .A1(n110), .A2(n334), .ZN(n53) );
  OR2_X1 U106 ( .A1(n416), .A2(n246), .ZN(n54) );
  NAND3_X1 U107 ( .A1(n54), .A2(n53), .A3(n176), .ZN(n225) );
  OR2_X1 U108 ( .A1(n25), .A2(n477), .ZN(n55) );
  OR2_X1 U109 ( .A1(n221), .A2(n246), .ZN(n56) );
  NAND3_X1 U110 ( .A1(n55), .A2(n56), .A3(n220), .ZN(n272) );
  OR2_X1 U111 ( .A1(n110), .A2(n463), .ZN(n57) );
  OR2_X1 U112 ( .A1(n210), .A2(n246), .ZN(n58) );
  NAND3_X1 U113 ( .A1(n57), .A2(n58), .A3(n209), .ZN(n262) );
  OR2_X1 U114 ( .A1(n37), .A2(n343), .ZN(n59) );
  OR2_X1 U115 ( .A1(n110), .A2(n425), .ZN(n60) );
  NAND3_X1 U116 ( .A1(n59), .A2(n60), .A3(n266), .ZN(n309) );
  MUX2_X1 U117 ( .A(n20), .B(n336), .S(n132), .Z(n326) );
  OR2_X1 U118 ( .A1(n25), .A2(n354), .ZN(n61) );
  OR2_X1 U119 ( .A1(n441), .A2(n246), .ZN(n62) );
  NAND3_X1 U120 ( .A1(n61), .A2(n62), .A3(n190), .ZN(n241) );
  OR2_X1 U121 ( .A1(n108), .A2(n477), .ZN(n63) );
  OR2_X1 U122 ( .A1(n110), .A2(n476), .ZN(n64) );
  NAND3_X1 U123 ( .A1(n63), .A2(n303), .A3(n64), .ZN(n349) );
  OR2_X1 U124 ( .A1(n452), .A2(n25), .ZN(n65) );
  OR2_X1 U125 ( .A1(n200), .A2(n246), .ZN(n66) );
  NAND3_X1 U126 ( .A1(n65), .A2(n66), .A3(n199), .ZN(n252) );
  OR2_X1 U127 ( .A1(n25), .A2(n343), .ZN(n67) );
  OR2_X1 U128 ( .A1(n428), .A2(n246), .ZN(n68) );
  NAND3_X1 U129 ( .A1(n67), .A2(n68), .A3(n185), .ZN(n231) );
  BUF_X1 U130 ( .A(n501), .Z(n107) );
  NAND2_X1 U131 ( .A1(DATA1[3]), .A2(n72), .ZN(n81) );
  INV_X1 U132 ( .A(n78), .ZN(n69) );
  OR2_X1 U133 ( .A1(n110), .A2(n405), .ZN(n70) );
  OR2_X1 U134 ( .A1(n502), .A2(n246), .ZN(n71) );
  NAND3_X1 U135 ( .A1(n245), .A2(n71), .A3(n70), .ZN(n291) );
  INV_X1 U136 ( .A(n107), .ZN(n72) );
  INV_X1 U137 ( .A(n107), .ZN(n474) );
  BUF_X2 U138 ( .A(n73), .Z(n110) );
  NAND3_X1 U139 ( .A1(n332), .A2(n103), .A3(n118), .ZN(n73) );
  OR2_X1 U140 ( .A1(n110), .A2(n441), .ZN(n74) );
  NAND2_X1 U141 ( .A1(n440), .A2(n74), .ZN(n489) );
  MUX2_X1 U142 ( .A(n356), .B(n76), .S(n140), .Z(n367) );
  INV_X1 U143 ( .A(n139), .ZN(n137) );
  MUX2_X1 U144 ( .A(n45), .B(n464), .S(n147), .Z(n417) );
  NOR2_X1 U145 ( .A1(n437), .A2(n10), .ZN(n439) );
  NAND3_X1 U146 ( .A1(n96), .A2(n97), .A3(n323), .ZN(n75) );
  INV_X1 U147 ( .A(n355), .ZN(n76) );
  MUX2_X1 U148 ( .A(n76), .B(n356), .S(n137), .Z(n77) );
  NAND3_X1 U149 ( .A1(n81), .A2(n82), .A3(n285), .ZN(n79) );
  BUF_X1 U150 ( .A(CONF), .Z(n117) );
  OR2_X1 U151 ( .A1(n25), .A2(n428), .ZN(n80) );
  NAND2_X1 U152 ( .A1(n80), .A2(n427), .ZN(n479) );
  OR2_X1 U153 ( .A1(n25), .A2(n451), .ZN(n82) );
  NAND3_X1 U154 ( .A1(n81), .A2(n82), .A3(n285), .ZN(n328) );
  BUF_X1 U155 ( .A(n478), .Z(n83) );
  OR2_X1 U156 ( .A1(n110), .A2(n416), .ZN(n84) );
  NAND2_X1 U157 ( .A1(n415), .A2(n84), .ZN(n464) );
  NAND2_X1 U158 ( .A1(n474), .A2(DATA1[16]), .ZN(n85) );
  NAND2_X1 U159 ( .A1(DATA1[0]), .A2(n505), .ZN(n86) );
  AND3_X1 U160 ( .A1(n85), .A2(n86), .A3(n9), .ZN(n415) );
  INV_X1 U161 ( .A(n11), .ZN(n87) );
  OR2_X1 U162 ( .A1(n37), .A2(n334), .ZN(n88) );
  OR2_X1 U163 ( .A1(n25), .A2(n414), .ZN(n89) );
  NAND3_X1 U164 ( .A1(n88), .A2(n89), .A3(n256), .ZN(n300) );
  INV_X1 U165 ( .A(n78), .ZN(n91) );
  INV_X1 U166 ( .A(n142), .ZN(n92) );
  AND2_X1 U167 ( .A1(n332), .A2(n126), .ZN(n93) );
  INV_X1 U168 ( .A(n160), .ZN(n94) );
  INV_X1 U169 ( .A(n160), .ZN(n95) );
  OR2_X1 U170 ( .A1(n108), .A2(n405), .ZN(n96) );
  OR2_X1 U171 ( .A1(n110), .A2(n404), .ZN(n97) );
  NAND3_X1 U172 ( .A1(n96), .A2(n97), .A3(n323), .ZN(n370) );
  INV_X1 U173 ( .A(n99), .ZN(n98) );
  INV_X1 U174 ( .A(DATA2[4]), .ZN(n99) );
  INV_X1 U175 ( .A(n103), .ZN(n100) );
  OAI221_X1 U176 ( .B1(n91), .B2(n405), .C1(n37), .C2(n404), .A(n403), .ZN(
        n102) );
  INV_X1 U177 ( .A(DATA2[4]), .ZN(n103) );
  OAI221_X1 U178 ( .B1(n452), .B2(n69), .C1(n451), .C2(n108), .A(n364), .ZN(
        n104) );
  MUX2_X1 U179 ( .A(n399), .B(n447), .S(n146), .Z(n394) );
  INV_X1 U180 ( .A(n146), .ZN(n144) );
  OR2_X1 U181 ( .A1(n37), .A2(n463), .ZN(n105) );
  OR2_X1 U182 ( .A1(n25), .A2(n462), .ZN(n106) );
  INV_X1 U183 ( .A(n160), .ZN(n322) );
  CLKBUF_X1 U184 ( .A(n116), .Z(n121) );
  NAND3_X1 U185 ( .A1(n103), .A2(n118), .A3(n101), .ZN(n501) );
  BUF_X2 U186 ( .A(n117), .Z(n125) );
  CLKBUF_X1 U187 ( .A(n117), .Z(n126) );
  CLKBUF_X1 U188 ( .A(n117), .Z(n124) );
  INV_X1 U189 ( .A(CONF), .ZN(n118) );
  INV_X1 U190 ( .A(CONF), .ZN(n120) );
  INV_X1 U191 ( .A(n146), .ZN(n142) );
  INV_X1 U192 ( .A(n146), .ZN(n141) );
  INV_X1 U193 ( .A(n132), .ZN(n129) );
  INV_X1 U194 ( .A(n132), .ZN(n127) );
  AND2_X1 U195 ( .A1(n126), .A2(n100), .ZN(n109) );
  AOI221_X1 U196 ( .B1(DATA1[6]), .B2(n41), .C1(DATA1[14]), .C2(n504), .A(n488), .ZN(n491) );
  OAI221_X1 U197 ( .B1(n108), .B2(n354), .C1(n110), .C2(n438), .A(n276), .ZN(
        n318) );
  BUF_X2 U198 ( .A(n90), .Z(n114) );
  OR2_X1 U199 ( .A1(n69), .A2(n343), .ZN(n111) );
  OR2_X1 U200 ( .A1(n37), .A2(n425), .ZN(n112) );
  INV_X1 U201 ( .A(DATA2[2]), .ZN(n146) );
  INV_X1 U202 ( .A(CONF), .ZN(n119) );
  INV_X1 U203 ( .A(DATA2[0]), .ZN(n132) );
  INV_X1 U204 ( .A(DATA2[0]), .ZN(n133) );
  INV_X1 U205 ( .A(DATA2[1]), .ZN(n139) );
  INV_X1 U206 ( .A(n146), .ZN(n145) );
  INV_X1 U207 ( .A(DATA2[3]), .ZN(n332) );
  INV_X1 U208 ( .A(n36), .ZN(n163) );
  NAND2_X1 U209 ( .A1(n109), .A2(n8), .ZN(n171) );
  INV_X1 U210 ( .A(n171), .ZN(n162) );
  INV_X1 U211 ( .A(DATA1[8]), .ZN(n414) );
  INV_X1 U212 ( .A(DATA1[0]), .ZN(n334) );
  OAI22_X1 U213 ( .A1(n414), .A2(n87), .B1(n334), .B2(n159), .ZN(n148) );
  INV_X1 U214 ( .A(DATA1[20]), .ZN(n150) );
  INV_X1 U215 ( .A(DATA1[28]), .ZN(n210) );
  AOI22_X1 U216 ( .A1(n113), .A2(DATA1[4]), .B1(n94), .B2(DATA1[12]), .ZN(n149) );
  OAI221_X1 U217 ( .B1(n150), .B2(n36), .C1(n210), .C2(n171), .A(n149), .ZN(
        n181) );
  INV_X1 U218 ( .A(n181), .ZN(n151) );
  MUX2_X1 U219 ( .A(n152), .B(n151), .S(n141), .Z(n158) );
  INV_X1 U220 ( .A(DATA1[18]), .ZN(n154) );
  INV_X1 U221 ( .A(DATA1[26]), .ZN(n441) );
  AOI22_X1 U222 ( .A1(n115), .A2(DATA1[2]), .B1(n95), .B2(DATA1[10]), .ZN(n153) );
  OAI221_X1 U223 ( .B1(n154), .B2(n36), .C1(n441), .C2(n171), .A(n153), .ZN(
        n156) );
  INV_X1 U224 ( .A(DATA1[22]), .ZN(n486) );
  INV_X1 U225 ( .A(DATA1[30]), .ZN(n487) );
  AOI22_X1 U226 ( .A1(n115), .A2(DATA1[6]), .B1(n95), .B2(DATA1[14]), .ZN(n155) );
  OAI221_X1 U227 ( .B1(n486), .B2(n36), .C1(n487), .C2(n171), .A(n155), .ZN(
        n203) );
  MUX2_X1 U228 ( .A(n156), .B(n203), .S(n141), .Z(n157) );
  INV_X1 U229 ( .A(n157), .ZN(n183) );
  MUX2_X1 U230 ( .A(n158), .B(n183), .S(n134), .Z(n175) );
  INV_X1 U231 ( .A(DATA1[9]), .ZN(n425) );
  INV_X1 U232 ( .A(DATA1[1]), .ZN(n343) );
  OAI22_X1 U233 ( .A1(n425), .A2(n87), .B1(n343), .B2(n159), .ZN(n161) );
  AOI221_X1 U234 ( .B1(n163), .B2(DATA1[17]), .C1(n162), .C2(DATA1[25]), .A(
        n161), .ZN(n167) );
  INV_X1 U235 ( .A(DATA1[21]), .ZN(n165) );
  INV_X1 U236 ( .A(DATA1[29]), .ZN(n221) );
  AOI22_X1 U237 ( .A1(n16), .A2(DATA1[5]), .B1(n11), .B2(DATA1[13]), .ZN(n164)
         );
  OAI221_X1 U238 ( .B1(n165), .B2(n36), .C1(n221), .C2(n171), .A(n164), .ZN(
        n193) );
  INV_X1 U239 ( .A(n193), .ZN(n166) );
  INV_X1 U240 ( .A(DATA1[19]), .ZN(n169) );
  INV_X1 U241 ( .A(DATA1[27]), .ZN(n200) );
  AOI22_X1 U242 ( .A1(n16), .A2(DATA1[3]), .B1(n94), .B2(DATA1[11]), .ZN(n168)
         );
  OAI221_X1 U243 ( .B1(n169), .B2(n36), .C1(n200), .C2(n171), .A(n168), .ZN(
        n172) );
  INV_X1 U244 ( .A(DATA1[23]), .ZN(n500) );
  INV_X1 U245 ( .A(DATA1[31]), .ZN(n502) );
  AOI22_X1 U246 ( .A1(n115), .A2(DATA1[7]), .B1(n95), .B2(DATA1[15]), .ZN(n170) );
  OAI221_X1 U247 ( .B1(n500), .B2(n36), .C1(n502), .C2(n171), .A(n170), .ZN(
        n214) );
  MUX2_X1 U248 ( .A(n172), .B(n214), .S(n141), .Z(n173) );
  INV_X1 U249 ( .A(n173), .ZN(n195) );
  MUX2_X1 U250 ( .A(n174), .B(n195), .S(n134), .Z(n184) );
  MUX2_X1 U251 ( .A(n175), .B(n184), .S(n127), .Z(n180) );
  INV_X1 U252 ( .A(DATA1[24]), .ZN(n416) );
  AOI22_X1 U253 ( .A1(n23), .A2(DATA1[8]), .B1(n95), .B2(DATA1[16]), .ZN(n176)
         );
  NAND2_X1 U254 ( .A1(n225), .A2(n147), .ZN(n191) );
  INV_X1 U255 ( .A(n191), .ZN(n177) );
  NAND2_X1 U256 ( .A1(n177), .A2(n140), .ZN(n187) );
  INV_X1 U257 ( .A(n187), .ZN(n178) );
  NAND3_X1 U258 ( .A1(n133), .A2(n178), .A3(n118), .ZN(n179) );
  NAND2_X1 U259 ( .A1(n180), .A2(n179), .ZN(OUTPUT[0]) );
  MUX2_X1 U260 ( .A(n181), .B(n225), .S(n141), .Z(n182) );
  INV_X1 U261 ( .A(n182), .ZN(n205) );
  MUX2_X1 U262 ( .A(n183), .B(n205), .S(n134), .Z(n196) );
  MUX2_X1 U263 ( .A(n184), .B(n196), .S(n127), .Z(n189) );
  INV_X1 U264 ( .A(DATA1[25]), .ZN(n428) );
  AOI22_X1 U265 ( .A1(n113), .A2(DATA1[9]), .B1(n94), .B2(DATA1[17]), .ZN(n185) );
  NAND2_X1 U266 ( .A1(n13), .A2(n147), .ZN(n201) );
  INV_X1 U267 ( .A(n201), .ZN(n186) );
  NAND2_X1 U268 ( .A1(n186), .A2(n140), .ZN(n192) );
  MUX2_X1 U269 ( .A(n192), .B(n187), .S(n127), .Z(n188) );
  OAI22_X1 U270 ( .A1(n189), .A2(n120), .B1(n125), .B2(n188), .ZN(OUTPUT[1])
         );
  INV_X1 U271 ( .A(DATA1[2]), .ZN(n354) );
  AOI22_X1 U272 ( .A1(n115), .A2(DATA1[10]), .B1(n11), .B2(DATA1[18]), .ZN(
        n190) );
  NAND2_X1 U273 ( .A1(n3), .A2(n147), .ZN(n212) );
  MUX2_X1 U274 ( .A(n212), .B(n191), .S(n134), .Z(n202) );
  MUX2_X1 U275 ( .A(n202), .B(n192), .S(n127), .Z(n198) );
  MUX2_X1 U276 ( .A(n193), .B(n231), .S(n141), .Z(n194) );
  INV_X1 U277 ( .A(n194), .ZN(n216) );
  MUX2_X1 U278 ( .A(n195), .B(n216), .S(n134), .Z(n206) );
  MUX2_X1 U279 ( .A(n196), .B(n206), .S(n127), .Z(n197) );
  OAI22_X1 U280 ( .A1(n121), .A2(n198), .B1(n197), .B2(n118), .ZN(OUTPUT[2])
         );
  INV_X1 U281 ( .A(DATA1[3]), .ZN(n452) );
  AOI22_X1 U282 ( .A1(n23), .A2(DATA1[11]), .B1(n94), .B2(DATA1[19]), .ZN(n199) );
  NAND2_X1 U283 ( .A1(n14), .A2(n147), .ZN(n223) );
  MUX2_X1 U284 ( .A(n223), .B(n201), .S(n134), .Z(n213) );
  MUX2_X1 U285 ( .A(n213), .B(n202), .S(n127), .Z(n208) );
  MUX2_X1 U286 ( .A(n203), .B(n241), .S(n141), .Z(n204) );
  INV_X1 U287 ( .A(n204), .ZN(n227) );
  MUX2_X1 U288 ( .A(n205), .B(n227), .S(n134), .Z(n217) );
  MUX2_X1 U289 ( .A(n206), .B(n217), .S(n127), .Z(n207) );
  OAI22_X1 U290 ( .A1(n121), .A2(n208), .B1(n207), .B2(n118), .ZN(OUTPUT[3])
         );
  INV_X1 U291 ( .A(DATA1[4]), .ZN(n463) );
  AOI22_X1 U292 ( .A1(n113), .A2(DATA1[12]), .B1(n94), .B2(DATA1[20]), .ZN(
        n209) );
  MUX2_X1 U293 ( .A(n262), .B(n225), .S(n141), .Z(n211) );
  INV_X1 U294 ( .A(n211), .ZN(n237) );
  MUX2_X1 U295 ( .A(n237), .B(n212), .S(n134), .Z(n224) );
  MUX2_X1 U296 ( .A(n224), .B(n213), .S(n127), .Z(n219) );
  MUX2_X1 U297 ( .A(n214), .B(n252), .S(n141), .Z(n215) );
  INV_X1 U298 ( .A(n215), .ZN(n233) );
  MUX2_X1 U299 ( .A(n217), .B(n228), .S(n127), .Z(n218) );
  OAI22_X1 U300 ( .A1(n121), .A2(n219), .B1(n218), .B2(n118), .ZN(OUTPUT[4])
         );
  INV_X1 U301 ( .A(DATA1[5]), .ZN(n477) );
  AOI22_X1 U302 ( .A1(n115), .A2(DATA1[13]), .B1(n11), .B2(DATA1[21]), .ZN(
        n220) );
  MUX2_X1 U303 ( .A(n272), .B(n13), .S(n141), .Z(n222) );
  INV_X1 U304 ( .A(n222), .ZN(n248) );
  MUX2_X1 U305 ( .A(n248), .B(n223), .S(n134), .Z(n238) );
  MUX2_X1 U306 ( .A(n238), .B(n224), .S(n127), .Z(n230) );
  MUX2_X1 U307 ( .A(n225), .B(n262), .S(n141), .Z(n226) );
  INV_X1 U308 ( .A(n226), .ZN(n243) );
  MUX2_X1 U309 ( .A(n227), .B(n243), .S(n134), .Z(n234) );
  MUX2_X1 U310 ( .A(n228), .B(n234), .S(n127), .Z(n229) );
  OAI22_X1 U311 ( .A1(n122), .A2(n230), .B1(n229), .B2(n118), .ZN(OUTPUT[5])
         );
  MUX2_X1 U312 ( .A(n231), .B(n272), .S(n141), .Z(n232) );
  INV_X1 U313 ( .A(n232), .ZN(n254) );
  MUX2_X1 U314 ( .A(n233), .B(n254), .S(n134), .Z(n244) );
  MUX2_X1 U315 ( .A(n234), .B(n244), .S(n127), .Z(n240) );
  INV_X1 U316 ( .A(DATA1[6]), .ZN(n393) );
  AOI22_X1 U317 ( .A1(n23), .A2(DATA1[14]), .B1(n95), .B2(DATA1[22]), .ZN(n235) );
  MUX2_X1 U318 ( .A(n42), .B(n241), .S(n142), .Z(n236) );
  INV_X1 U319 ( .A(n236), .ZN(n258) );
  MUX2_X1 U320 ( .A(n258), .B(n237), .S(n135), .Z(n249) );
  MUX2_X1 U321 ( .A(n249), .B(n238), .S(n128), .Z(n239) );
  OAI22_X1 U322 ( .A1(n240), .A2(n119), .B1(n239), .B2(n125), .ZN(OUTPUT[6])
         );
  MUX2_X1 U323 ( .A(n3), .B(n42), .S(n142), .Z(n242) );
  INV_X1 U324 ( .A(n242), .ZN(n264) );
  MUX2_X1 U325 ( .A(n243), .B(n264), .S(n135), .Z(n255) );
  MUX2_X1 U326 ( .A(n244), .B(n255), .S(n128), .Z(n251) );
  INV_X1 U327 ( .A(DATA1[7]), .ZN(n405) );
  AOI22_X1 U328 ( .A1(n115), .A2(DATA1[15]), .B1(n95), .B2(DATA1[23]), .ZN(
        n245) );
  INV_X1 U329 ( .A(n247), .ZN(n268) );
  MUX2_X1 U330 ( .A(n268), .B(n248), .S(n135), .Z(n259) );
  OAI22_X1 U331 ( .A1(n251), .A2(n118), .B1(n250), .B2(n125), .ZN(OUTPUT[7])
         );
  MUX2_X1 U332 ( .A(n252), .B(n291), .S(n142), .Z(n253) );
  INV_X1 U333 ( .A(n253), .ZN(n274) );
  MUX2_X1 U334 ( .A(n254), .B(n274), .S(n135), .Z(n265) );
  MUX2_X1 U335 ( .A(n255), .B(n265), .S(n128), .Z(n261) );
  AOI22_X1 U336 ( .A1(n23), .A2(DATA1[16]), .B1(n11), .B2(DATA1[24]), .ZN(n256) );
  MUX2_X1 U337 ( .A(n300), .B(n262), .S(n142), .Z(n257) );
  INV_X1 U338 ( .A(n257), .ZN(n278) );
  MUX2_X1 U339 ( .A(n278), .B(n258), .S(n135), .Z(n269) );
  MUX2_X1 U340 ( .A(n269), .B(n259), .S(n128), .Z(n260) );
  OAI22_X1 U341 ( .A1(n261), .A2(n119), .B1(n260), .B2(n125), .ZN(OUTPUT[8])
         );
  MUX2_X1 U342 ( .A(n262), .B(n18), .S(n142), .Z(n263) );
  INV_X1 U343 ( .A(n263), .ZN(n283) );
  MUX2_X1 U344 ( .A(n264), .B(n283), .S(n135), .Z(n275) );
  MUX2_X1 U345 ( .A(n265), .B(n275), .S(n128), .Z(n271) );
  AOI22_X1 U346 ( .A1(n16), .A2(DATA1[17]), .B1(n11), .B2(DATA1[25]), .ZN(n266) );
  MUX2_X1 U347 ( .A(n309), .B(n272), .S(n142), .Z(n267) );
  INV_X1 U348 ( .A(n267), .ZN(n287) );
  MUX2_X1 U349 ( .A(n287), .B(n268), .S(n135), .Z(n279) );
  MUX2_X1 U350 ( .A(n279), .B(n269), .S(n128), .Z(n270) );
  OAI22_X1 U351 ( .A1(n271), .A2(n119), .B1(n270), .B2(n125), .ZN(OUTPUT[9])
         );
  MUX2_X1 U352 ( .A(n272), .B(n17), .S(n142), .Z(n273) );
  INV_X1 U353 ( .A(n273), .ZN(n292) );
  MUX2_X1 U354 ( .A(n274), .B(n292), .S(n135), .Z(n284) );
  MUX2_X1 U355 ( .A(n275), .B(n284), .S(n128), .Z(n281) );
  INV_X1 U356 ( .A(DATA1[10]), .ZN(n438) );
  AOI22_X1 U357 ( .A1(n114), .A2(DATA1[18]), .B1(n322), .B2(DATA1[26]), .ZN(
        n276) );
  INV_X1 U358 ( .A(n277), .ZN(n296) );
  MUX2_X1 U359 ( .A(n288), .B(n279), .S(n128), .Z(n280) );
  OAI22_X1 U360 ( .A1(n281), .A2(n119), .B1(n280), .B2(n124), .ZN(OUTPUT[10])
         );
  MUX2_X1 U361 ( .A(n42), .B(n318), .S(n142), .Z(n282) );
  MUX2_X1 U362 ( .A(n283), .B(n21), .S(n135), .Z(n293) );
  MUX2_X1 U363 ( .A(n284), .B(n293), .S(n128), .Z(n290) );
  INV_X1 U364 ( .A(DATA1[11]), .ZN(n451) );
  AOI22_X1 U365 ( .A1(n115), .A2(DATA1[19]), .B1(n94), .B2(DATA1[27]), .ZN(
        n285) );
  INV_X1 U366 ( .A(n286), .ZN(n305) );
  MUX2_X1 U367 ( .A(n305), .B(n287), .S(n135), .Z(n297) );
  MUX2_X1 U368 ( .A(n297), .B(n288), .S(n128), .Z(n289) );
  OAI22_X1 U369 ( .A1(n290), .A2(n119), .B1(n289), .B2(n124), .ZN(OUTPUT[11])
         );
  MUX2_X1 U370 ( .A(n292), .B(n38), .S(n135), .Z(n302) );
  MUX2_X1 U371 ( .A(n293), .B(n302), .S(n128), .Z(n299) );
  INV_X1 U372 ( .A(DATA1[12]), .ZN(n462) );
  AOI22_X1 U373 ( .A1(n115), .A2(DATA1[20]), .B1(n322), .B2(DATA1[28]), .ZN(
        n294) );
  INV_X1 U374 ( .A(n295), .ZN(n314) );
  MUX2_X1 U375 ( .A(n314), .B(n296), .S(n136), .Z(n306) );
  MUX2_X1 U376 ( .A(n306), .B(n297), .S(n129), .Z(n298) );
  OAI22_X1 U377 ( .A1(n299), .A2(n119), .B1(n298), .B2(n124), .ZN(OUTPUT[12])
         );
  MUX2_X1 U378 ( .A(n300), .B(n19), .S(n143), .Z(n301) );
  INV_X1 U379 ( .A(n301), .ZN(n320) );
  MUX2_X1 U380 ( .A(n21), .B(n320), .S(n136), .Z(n311) );
  MUX2_X1 U381 ( .A(n302), .B(n311), .S(n129), .Z(n308) );
  INV_X1 U382 ( .A(DATA1[13]), .ZN(n476) );
  AOI22_X1 U383 ( .A1(n115), .A2(DATA1[21]), .B1(n322), .B2(DATA1[29]), .ZN(
        n303) );
  MUX2_X1 U384 ( .A(n349), .B(n309), .S(n143), .Z(n304) );
  INV_X1 U385 ( .A(n304), .ZN(n325) );
  MUX2_X1 U386 ( .A(n315), .B(n306), .S(n129), .Z(n307) );
  OAI22_X1 U387 ( .A1(n308), .A2(n119), .B1(n307), .B2(n124), .ZN(OUTPUT[13])
         );
  MUX2_X1 U388 ( .A(n17), .B(n349), .S(n143), .Z(n310) );
  INV_X1 U389 ( .A(n310), .ZN(n330) );
  MUX2_X1 U390 ( .A(n311), .B(n321), .S(n129), .Z(n317) );
  INV_X1 U391 ( .A(DATA1[14]), .ZN(n392) );
  AOI22_X1 U392 ( .A1(n113), .A2(DATA1[22]), .B1(n322), .B2(DATA1[30]), .ZN(
        n312) );
  MUX2_X1 U393 ( .A(n360), .B(n318), .S(n143), .Z(n313) );
  MUX2_X1 U394 ( .A(n20), .B(n315), .S(n129), .Z(n316) );
  OAI22_X1 U395 ( .A1(n317), .A2(n119), .B1(n316), .B2(n124), .ZN(OUTPUT[14])
         );
  MUX2_X1 U396 ( .A(n318), .B(n360), .S(n143), .Z(n319) );
  INV_X1 U397 ( .A(n319), .ZN(n340) );
  MUX2_X1 U398 ( .A(n320), .B(n340), .S(n136), .Z(n331) );
  MUX2_X1 U399 ( .A(n321), .B(n331), .S(n129), .Z(n327) );
  INV_X1 U400 ( .A(DATA1[15]), .ZN(n404) );
  AOI22_X1 U401 ( .A1(n16), .A2(DATA1[23]), .B1(n322), .B2(DATA1[31]), .ZN(
        n323) );
  MUX2_X1 U402 ( .A(n370), .B(n328), .S(n143), .Z(n324) );
  INV_X1 U403 ( .A(n324), .ZN(n345) );
  MUX2_X1 U404 ( .A(n345), .B(n325), .S(n136), .Z(n336) );
  OAI22_X1 U405 ( .A1(n327), .A2(n119), .B1(n326), .B2(n124), .ZN(OUTPUT[15])
         );
  MUX2_X1 U406 ( .A(n79), .B(n75), .S(n143), .Z(n329) );
  INV_X1 U407 ( .A(n329), .ZN(n351) );
  MUX2_X1 U408 ( .A(n330), .B(n351), .S(n136), .Z(n341) );
  MUX2_X1 U409 ( .A(n331), .B(n341), .S(n129), .Z(n338) );
  AOI22_X1 U410 ( .A1(n27), .A2(DATA1[16]), .B1(n114), .B2(DATA1[24]), .ZN(
        n333) );
  MUX2_X1 U411 ( .A(n379), .B(n19), .S(n143), .Z(n335) );
  INV_X1 U412 ( .A(n335), .ZN(n356) );
  MUX2_X1 U413 ( .A(n356), .B(n22), .S(n136), .Z(n346) );
  OAI22_X1 U414 ( .A1(n338), .A2(n119), .B1(n337), .B2(n123), .ZN(OUTPUT[16])
         );
  MUX2_X1 U415 ( .A(n19), .B(n379), .S(n143), .Z(n339) );
  INV_X1 U416 ( .A(n339), .ZN(n362) );
  MUX2_X1 U417 ( .A(n340), .B(n362), .S(n136), .Z(n352) );
  MUX2_X1 U418 ( .A(n341), .B(n352), .S(n129), .Z(n348) );
  AOI22_X1 U419 ( .A1(DATA1[17]), .A2(n27), .B1(n115), .B2(DATA1[25]), .ZN(
        n342) );
  MUX2_X1 U420 ( .A(n46), .B(n349), .S(n143), .Z(n344) );
  INV_X1 U421 ( .A(n344), .ZN(n366) );
  MUX2_X1 U422 ( .A(n366), .B(n345), .S(n136), .Z(n357) );
  MUX2_X1 U423 ( .A(n357), .B(n32), .S(n129), .Z(n347) );
  OAI22_X1 U424 ( .A1(n348), .A2(n119), .B1(n347), .B2(n123), .ZN(OUTPUT[17])
         );
  MUX2_X1 U425 ( .A(n349), .B(n46), .S(n143), .Z(n350) );
  INV_X1 U426 ( .A(n350), .ZN(n372) );
  MUX2_X1 U427 ( .A(n351), .B(n372), .S(n136), .Z(n363) );
  MUX2_X1 U428 ( .A(n352), .B(n363), .S(n129), .Z(n359) );
  AOI22_X1 U429 ( .A1(DATA1[18]), .A2(n27), .B1(n114), .B2(DATA1[26]), .ZN(
        n353) );
  OAI221_X1 U430 ( .B1(n69), .B2(n354), .C1(n108), .C2(n438), .A(n353), .ZN(
        n399) );
  MUX2_X1 U431 ( .A(n399), .B(n31), .S(n144), .Z(n355) );
  MUX2_X1 U432 ( .A(n77), .B(n357), .S(n130), .Z(n358) );
  OAI22_X1 U433 ( .A1(n359), .A2(n120), .B1(n358), .B2(n123), .ZN(OUTPUT[18])
         );
  MUX2_X1 U434 ( .A(n31), .B(n399), .S(n144), .Z(n361) );
  INV_X1 U435 ( .A(n361), .ZN(n381) );
  MUX2_X1 U436 ( .A(n362), .B(n381), .S(n137), .Z(n373) );
  MUX2_X1 U437 ( .A(n363), .B(n373), .S(n130), .Z(n369) );
  AOI22_X1 U438 ( .A1(n27), .A2(DATA1[19]), .B1(n114), .B2(DATA1[27]), .ZN(
        n364) );
  MUX2_X1 U439 ( .A(n104), .B(n370), .S(n144), .Z(n365) );
  INV_X1 U440 ( .A(n365), .ZN(n385) );
  MUX2_X1 U441 ( .A(n385), .B(n366), .S(n137), .Z(n376) );
  MUX2_X1 U442 ( .A(n376), .B(n367), .S(n130), .Z(n368) );
  OAI22_X1 U443 ( .A1(n369), .A2(n119), .B1(n368), .B2(n123), .ZN(OUTPUT[19])
         );
  MUX2_X1 U444 ( .A(n75), .B(n104), .S(n144), .Z(n371) );
  INV_X1 U445 ( .A(n371), .ZN(n389) );
  MUX2_X1 U446 ( .A(n372), .B(n389), .S(n137), .Z(n382) );
  MUX2_X1 U447 ( .A(n373), .B(n382), .S(n130), .Z(n378) );
  AOI22_X1 U448 ( .A1(DATA1[20]), .A2(n27), .B1(n114), .B2(DATA1[28]), .ZN(
        n374) );
  MUX2_X1 U449 ( .A(n422), .B(n379), .S(n144), .Z(n375) );
  INV_X1 U450 ( .A(n375), .ZN(n395) );
  MUX2_X1 U451 ( .A(n30), .B(n376), .S(n130), .Z(n377) );
  OAI22_X1 U452 ( .A1(n378), .A2(n120), .B1(n377), .B2(n123), .ZN(OUTPUT[20])
         );
  MUX2_X1 U453 ( .A(n379), .B(n422), .S(n144), .Z(n380) );
  INV_X1 U454 ( .A(n380), .ZN(n401) );
  MUX2_X1 U455 ( .A(n381), .B(n401), .S(n137), .Z(n390) );
  MUX2_X1 U456 ( .A(n382), .B(n390), .S(n130), .Z(n387) );
  AOI22_X1 U457 ( .A1(DATA1[21]), .A2(n27), .B1(n23), .B2(DATA1[29]), .ZN(n383) );
  INV_X1 U458 ( .A(n384), .ZN(n407) );
  MUX2_X1 U459 ( .A(n407), .B(n385), .S(n137), .Z(n396) );
  MUX2_X1 U460 ( .A(n396), .B(n30), .S(n130), .Z(n386) );
  OAI22_X1 U461 ( .A1(n387), .A2(n120), .B1(n386), .B2(n123), .ZN(OUTPUT[21])
         );
  MUX2_X1 U462 ( .A(n1), .B(n434), .S(n144), .Z(n388) );
  INV_X1 U463 ( .A(n388), .ZN(n412) );
  MUX2_X1 U464 ( .A(n389), .B(n412), .S(n137), .Z(n402) );
  MUX2_X1 U465 ( .A(n390), .B(n402), .S(n130), .Z(n398) );
  AOI22_X1 U466 ( .A1(DATA1[22]), .A2(n27), .B1(n115), .B2(DATA1[30]), .ZN(
        n391) );
  INV_X1 U467 ( .A(n394), .ZN(n418) );
  MUX2_X1 U468 ( .A(n408), .B(n396), .S(n130), .Z(n397) );
  OAI22_X1 U469 ( .A1(n398), .A2(n120), .B1(n123), .B2(n397), .ZN(OUTPUT[22])
         );
  MUX2_X1 U470 ( .A(n399), .B(n447), .S(n144), .Z(n400) );
  INV_X1 U471 ( .A(n400), .ZN(n423) );
  MUX2_X1 U472 ( .A(n401), .B(n423), .S(n137), .Z(n413) );
  MUX2_X1 U473 ( .A(n402), .B(n413), .S(n130), .Z(n410) );
  OAI221_X1 U474 ( .B1(n91), .B2(n405), .C1(n108), .C2(n404), .A(n403), .ZN(
        n458) );
  INV_X1 U475 ( .A(n406), .ZN(n430) );
  MUX2_X1 U476 ( .A(n419), .B(n408), .S(n130), .Z(n409) );
  OAI22_X1 U477 ( .A1(n410), .A2(n120), .B1(n409), .B2(n124), .ZN(OUTPUT[23])
         );
  MUX2_X1 U478 ( .A(n104), .B(n458), .S(n144), .Z(n411) );
  INV_X1 U479 ( .A(n411), .ZN(n435) );
  MUX2_X1 U480 ( .A(n412), .B(n435), .S(n137), .Z(n424) );
  MUX2_X1 U481 ( .A(n413), .B(n424), .S(n130), .Z(n421) );
  NAND3_X1 U482 ( .A1(n8), .A2(n100), .A3(n118), .ZN(n478) );
  INV_X1 U483 ( .A(n478), .ZN(n505) );
  NAND2_X1 U484 ( .A1(n98), .A2(n118), .ZN(n437) );
  INV_X1 U485 ( .A(n417), .ZN(n443) );
  MUX2_X1 U486 ( .A(n431), .B(n419), .S(n131), .Z(n420) );
  OAI22_X1 U487 ( .A1(n421), .A2(n120), .B1(n420), .B2(n122), .ZN(OUTPUT[24])
         );
  NAND2_X1 U488 ( .A1(n45), .A2(n147), .ZN(n448) );
  MUX2_X1 U489 ( .A(n423), .B(n448), .S(n138), .Z(n436) );
  MUX2_X1 U490 ( .A(n424), .B(n436), .S(n131), .Z(n433) );
  NOR3_X1 U491 ( .A1(n425), .A2(n8), .A3(n437), .ZN(n426) );
  AOI221_X1 U492 ( .B1(n474), .B2(DATA1[17]), .C1(DATA1[1]), .C2(n41), .A(n426), .ZN(n427) );
  MUX2_X1 U493 ( .A(n479), .B(n33), .S(n145), .Z(n429) );
  INV_X1 U494 ( .A(n429), .ZN(n454) );
  OAI22_X1 U495 ( .A1(n433), .A2(n120), .B1(n432), .B2(n122), .ZN(OUTPUT[25])
         );
  NAND2_X1 U496 ( .A1(n33), .A2(n147), .ZN(n459) );
  MUX2_X1 U497 ( .A(n435), .B(n459), .S(n138), .Z(n449) );
  MUX2_X1 U498 ( .A(n436), .B(n449), .S(n131), .Z(n446) );
  AOI221_X1 U499 ( .B1(n474), .B2(DATA1[18]), .C1(DATA1[2]), .C2(n505), .A(
        n439), .ZN(n440) );
  MUX2_X1 U500 ( .A(n489), .B(n12), .S(n145), .Z(n442) );
  INV_X1 U501 ( .A(n442), .ZN(n467) );
  MUX2_X1 U502 ( .A(n455), .B(n444), .S(n131), .Z(n445) );
  OAI22_X1 U503 ( .A1(n446), .A2(n120), .B1(n445), .B2(n122), .ZN(OUTPUT[26])
         );
  NAND2_X1 U504 ( .A1(n12), .A2(n147), .ZN(n471) );
  MUX2_X1 U505 ( .A(n448), .B(n471), .S(n138), .Z(n460) );
  MUX2_X1 U506 ( .A(n449), .B(n460), .S(n131), .Z(n457) );
  AOI22_X1 U507 ( .A1(DATA1[19]), .A2(n72), .B1(n27), .B2(DATA1[27]), .ZN(n450) );
  MUX2_X1 U508 ( .A(n506), .B(n102), .S(n145), .Z(n453) );
  INV_X1 U509 ( .A(n453), .ZN(n482) );
  MUX2_X1 U510 ( .A(n482), .B(n454), .S(n138), .Z(n468) );
  MUX2_X1 U511 ( .A(n468), .B(n455), .S(n131), .Z(n456) );
  OAI22_X1 U512 ( .A1(n457), .A2(n120), .B1(n122), .B2(n456), .ZN(OUTPUT[27])
         );
  NAND2_X1 U513 ( .A1(n102), .A2(n147), .ZN(n495) );
  MUX2_X1 U514 ( .A(n459), .B(n495), .S(n138), .Z(n473) );
  MUX2_X1 U515 ( .A(n460), .B(n473), .S(n131), .Z(n470) );
  AOI22_X1 U516 ( .A1(DATA1[20]), .A2(n72), .B1(n27), .B2(DATA1[28]), .ZN(n461) );
  OAI221_X1 U517 ( .B1(n83), .B2(n463), .C1(n91), .C2(n462), .A(n461), .ZN(
        n465) );
  MUX2_X1 U518 ( .A(n465), .B(n464), .S(n145), .Z(n466) );
  INV_X1 U519 ( .A(n466), .ZN(n492) );
  MUX2_X1 U520 ( .A(n492), .B(n467), .S(n138), .Z(n483) );
  MUX2_X1 U521 ( .A(n483), .B(n468), .S(n131), .Z(n469) );
  OAI22_X1 U522 ( .A1(n470), .A2(n120), .B1(n469), .B2(n122), .ZN(OUTPUT[28])
         );
  INV_X1 U523 ( .A(n471), .ZN(n472) );
  NAND2_X1 U524 ( .A1(n472), .A2(n140), .ZN(n497) );
  MUX2_X1 U525 ( .A(n473), .B(n497), .S(n131), .Z(n485) );
  AOI22_X1 U526 ( .A1(DATA1[21]), .A2(n72), .B1(n2), .B2(DATA1[29]), .ZN(n475)
         );
  OAI221_X1 U527 ( .B1(n83), .B2(n477), .C1(n91), .C2(n476), .A(n475), .ZN(
        n480) );
  MUX2_X1 U528 ( .A(n480), .B(n479), .S(n145), .Z(n481) );
  INV_X1 U529 ( .A(n481), .ZN(n509) );
  MUX2_X1 U530 ( .A(n494), .B(n483), .S(n131), .Z(n484) );
  OAI22_X1 U531 ( .A1(n485), .A2(n120), .B1(n484), .B2(n122), .ZN(OUTPUT[29])
         );
  INV_X1 U532 ( .A(n69), .ZN(n504) );
  OAI22_X1 U533 ( .A1(n487), .A2(n110), .B1(n108), .B2(n486), .ZN(n488) );
  INV_X1 U534 ( .A(n489), .ZN(n490) );
  MUX2_X1 U535 ( .A(n491), .B(n490), .S(n145), .Z(n493) );
  MUX2_X1 U536 ( .A(n493), .B(n492), .S(n138), .Z(n511) );
  MUX2_X1 U537 ( .A(n511), .B(n494), .S(n131), .Z(n499) );
  INV_X1 U538 ( .A(n495), .ZN(n496) );
  NAND2_X1 U539 ( .A1(n496), .A2(n140), .ZN(n513) );
  MUX2_X1 U540 ( .A(n497), .B(n513), .S(n131), .Z(n498) );
  OAI22_X1 U541 ( .A1(n499), .A2(n121), .B1(n498), .B2(n118), .ZN(OUTPUT[30])
         );
  OAI22_X1 U542 ( .A1(n502), .A2(n25), .B1(n37), .B2(n500), .ZN(n503) );
  INV_X1 U543 ( .A(n34), .ZN(n507) );
  MUX2_X1 U544 ( .A(n508), .B(n507), .S(n145), .Z(n510) );
  MUX2_X1 U545 ( .A(n510), .B(n509), .S(n138), .Z(n512) );
  MUX2_X1 U546 ( .A(n512), .B(n511), .S(n130), .Z(n516) );
  INV_X1 U547 ( .A(n513), .ZN(n514) );
  NAND3_X1 U548 ( .A1(n133), .A2(n514), .A3(n125), .ZN(n515) );
  NAND2_X1 U549 ( .A1(n516), .A2(n515), .ZN(OUTPUT[31]) );
endmodule


module ALU_N32_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371;

  CLKBUF_X1 U3 ( .A(A[6]), .Z(n1) );
  XNOR2_X1 U4 ( .A(n124), .B(n2), .ZN(DIFF[30]) );
  NAND2_X1 U5 ( .A1(n123), .A2(n117), .ZN(n2) );
  NAND4_X1 U6 ( .A1(n206), .A2(n201), .A3(n202), .A4(n195), .ZN(n3) );
  AND2_X1 U7 ( .A1(n306), .A2(n280), .ZN(n4) );
  OR2_X1 U8 ( .A1(n339), .A2(A[12]), .ZN(n306) );
  AND2_X1 U9 ( .A1(n43), .A2(n9), .ZN(n5) );
  AND2_X1 U10 ( .A1(n169), .A2(n5), .ZN(n44) );
  CLKBUF_X1 U11 ( .A(A[10]), .Z(n6) );
  NAND3_X1 U12 ( .A1(n319), .A2(n318), .A3(n4), .ZN(n317) );
  BUF_X1 U13 ( .A(n325), .Z(n7) );
  CLKBUF_X1 U14 ( .A(n288), .Z(n8) );
  OAI21_X1 U15 ( .B1(n41), .B2(n295), .A(n89), .ZN(n76) );
  AND4_X1 U16 ( .A1(n306), .A2(n280), .A3(n282), .A4(n38), .ZN(n51) );
  AND2_X1 U17 ( .A1(n97), .A2(n29), .ZN(n18) );
  NAND2_X1 U18 ( .A1(n316), .A2(n280), .ZN(n315) );
  INV_X1 U19 ( .A(n18), .ZN(n95) );
  INV_X1 U20 ( .A(n36), .ZN(n154) );
  AND2_X1 U21 ( .A1(n160), .A2(n152), .ZN(n9) );
  AND2_X1 U22 ( .A1(n226), .A2(n206), .ZN(n10) );
  AND2_X1 U23 ( .A1(n76), .A2(n335), .ZN(n11) );
  AND2_X1 U24 ( .A1(n346), .A2(n72), .ZN(n12) );
  INV_X1 U25 ( .A(n82), .ZN(n13) );
  AND2_X1 U26 ( .A1(n114), .A2(n23), .ZN(n33) );
  AOI21_X1 U27 ( .B1(n352), .B2(n353), .A(n22), .ZN(n14) );
  CLKBUF_X1 U28 ( .A(n71), .Z(n15) );
  BUF_X1 U29 ( .A(n87), .Z(n16) );
  NAND2_X1 U30 ( .A1(n25), .A2(n10), .ZN(n17) );
  CLKBUF_X1 U31 ( .A(n111), .Z(n19) );
  AND2_X1 U32 ( .A1(n258), .A2(n257), .ZN(n20) );
  INV_X1 U33 ( .A(n283), .ZN(n21) );
  AND2_X1 U34 ( .A1(n354), .A2(n105), .ZN(n22) );
  AND2_X1 U35 ( .A1(n112), .A2(n113), .ZN(n23) );
  NOR2_X1 U36 ( .A1(n285), .A2(n27), .ZN(n24) );
  NAND2_X1 U37 ( .A1(n24), .A2(n273), .ZN(n25) );
  OR2_X1 U38 ( .A1(n344), .A2(A[11]), .ZN(n286) );
  XNOR2_X1 U39 ( .A(n309), .B(n26), .ZN(DIFF[14]) );
  AND2_X1 U40 ( .A1(n282), .A2(n278), .ZN(n26) );
  AND4_X1 U41 ( .A1(n297), .A2(n51), .A3(n283), .A4(n56), .ZN(n27) );
  NAND2_X1 U42 ( .A1(n77), .A2(n11), .ZN(n349) );
  NOR2_X1 U43 ( .A1(n27), .A2(n285), .ZN(n28) );
  NAND2_X1 U44 ( .A1(A[4]), .A2(n364), .ZN(n29) );
  NAND2_X1 U45 ( .A1(n201), .A2(n202), .ZN(n30) );
  NAND2_X1 U46 ( .A1(n216), .A2(n31), .ZN(n215) );
  INV_X1 U47 ( .A(n30), .ZN(n31) );
  NOR2_X1 U48 ( .A1(n65), .A2(A[0]), .ZN(n49) );
  CLKBUF_X1 U49 ( .A(n158), .Z(n32) );
  AND4_X1 U50 ( .A1(n99), .A2(n94), .A3(n87), .A4(n89), .ZN(n56) );
  XOR2_X1 U51 ( .A(n34), .B(n136), .Z(DIFF[29]) );
  AND2_X1 U52 ( .A1(n118), .A2(n122), .ZN(n34) );
  NOR2_X1 U53 ( .A1(n55), .A2(n49), .ZN(n35) );
  AND2_X1 U54 ( .A1(A[24]), .A2(n208), .ZN(n36) );
  NAND2_X1 U55 ( .A1(n14), .A2(n284), .ZN(n37) );
  NAND2_X1 U56 ( .A1(n14), .A2(n284), .ZN(n81) );
  NAND2_X1 U57 ( .A1(B[15]), .A2(n311), .ZN(n38) );
  NOR2_X1 U58 ( .A1(n231), .A2(n230), .ZN(n39) );
  NOR2_X1 U59 ( .A1(n39), .A2(n40), .ZN(n47) );
  OR2_X1 U60 ( .A1(n217), .A2(n229), .ZN(n40) );
  AND2_X1 U61 ( .A1(n362), .A2(n363), .ZN(n41) );
  NAND2_X1 U62 ( .A1(B[13]), .A2(n327), .ZN(n280) );
  NAND2_X1 U63 ( .A1(n28), .A2(n273), .ZN(n42) );
  NAND2_X1 U64 ( .A1(n272), .A2(n273), .ZN(n169) );
  NOR2_X1 U65 ( .A1(n227), .A2(n3), .ZN(n43) );
  NAND2_X1 U66 ( .A1(n17), .A2(n47), .ZN(n45) );
  AND2_X1 U67 ( .A1(n45), .A2(n46), .ZN(n218) );
  OR2_X1 U68 ( .A1(n217), .A2(n201), .ZN(n46) );
  CLKBUF_X1 U69 ( .A(A[5]), .Z(n48) );
  CLKBUF_X1 U70 ( .A(B[2]), .Z(n50) );
  AND3_X1 U71 ( .A1(n35), .A2(n105), .A3(n350), .ZN(n52) );
  AND2_X1 U72 ( .A1(n193), .A2(n53), .ZN(n273) );
  AND2_X1 U73 ( .A1(n192), .A2(n191), .ZN(n53) );
  XOR2_X1 U74 ( .A(n54), .B(n172), .Z(DIFF[26]) );
  AND2_X1 U75 ( .A1(n153), .A2(n158), .ZN(n54) );
  AND2_X1 U76 ( .A1(n317), .A2(n60), .ZN(n309) );
  AOI21_X1 U77 ( .B1(n133), .B2(n249), .A(n55), .ZN(n352) );
  OAI21_X1 U78 ( .B1(n78), .B2(n21), .A(n7), .ZN(n329) );
  NAND2_X1 U79 ( .A1(n21), .A2(n325), .ZN(n318) );
  NAND2_X1 U80 ( .A1(n323), .A2(n324), .ZN(n319) );
  AND2_X1 U81 ( .A1(n325), .A2(n76), .ZN(n323) );
  NAND2_X1 U82 ( .A1(n234), .A2(n231), .ZN(n233) );
  NAND2_X1 U83 ( .A1(n110), .A2(n111), .ZN(n109) );
  NOR2_X1 U84 ( .A1(n119), .A2(n59), .ZN(n108) );
  NOR2_X1 U85 ( .A1(n115), .A2(n116), .ZN(n110) );
  AND2_X1 U86 ( .A1(n66), .A2(n304), .ZN(n55) );
  NAND2_X1 U87 ( .A1(n175), .A2(n9), .ZN(n170) );
  NAND2_X1 U88 ( .A1(n49), .A2(n249), .ZN(n134) );
  NAND4_X1 U89 ( .A1(n334), .A2(n286), .A3(n71), .A4(n74), .ZN(n296) );
  XOR2_X1 U90 ( .A(n57), .B(n101), .Z(DIFF[3]) );
  AND2_X1 U91 ( .A1(n105), .A2(n106), .ZN(n57) );
  NAND2_X1 U92 ( .A1(n306), .A2(n277), .ZN(n328) );
  XNOR2_X1 U93 ( .A(n343), .B(n345), .ZN(DIFF[10]) );
  NAND4_X1 U94 ( .A1(n306), .A2(n280), .A3(n282), .A4(n281), .ZN(n289) );
  OAI21_X1 U95 ( .B1(n18), .B2(n92), .A(n93), .ZN(n88) );
  XNOR2_X1 U96 ( .A(n83), .B(n84), .ZN(DIFF[7]) );
  XOR2_X1 U97 ( .A(n69), .B(n70), .Z(DIFF[9]) );
  XNOR2_X1 U98 ( .A(n96), .B(n95), .ZN(DIFF[5]) );
  NAND2_X1 U99 ( .A1(n94), .A2(n93), .ZN(n96) );
  XNOR2_X1 U100 ( .A(n248), .B(n134), .ZN(DIFF[1]) );
  NAND2_X1 U101 ( .A1(n152), .A2(n159), .ZN(n179) );
  NAND2_X1 U102 ( .A1(n201), .A2(n199), .ZN(n222) );
  XNOR2_X1 U103 ( .A(n232), .B(n233), .ZN(DIFF[20]) );
  NAND2_X1 U104 ( .A1(n206), .A2(n200), .ZN(n232) );
  XNOR2_X1 U105 ( .A(n256), .B(n253), .ZN(DIFF[18]) );
  NAND2_X1 U106 ( .A1(n16), .A2(n85), .ZN(n91) );
  XNOR2_X1 U107 ( .A(n320), .B(n321), .ZN(DIFF[13]) );
  NAND2_X1 U108 ( .A1(n280), .A2(n279), .ZN(n320) );
  XNOR2_X1 U109 ( .A(n266), .B(n267), .ZN(DIFF[17]) );
  NAND2_X1 U110 ( .A1(n269), .A2(n262), .ZN(n266) );
  XNOR2_X1 U111 ( .A(n78), .B(n79), .ZN(DIFF[8]) );
  AOI21_X1 U112 ( .B1(n73), .B2(n74), .A(n75), .ZN(n69) );
  NAND2_X1 U113 ( .A1(n13), .A2(n77), .ZN(n73) );
  NAND2_X1 U114 ( .A1(n142), .A2(n141), .ZN(n149) );
  OAI21_X1 U115 ( .B1(n127), .B2(n120), .A(n118), .ZN(n126) );
  INV_X1 U116 ( .A(n63), .ZN(n350) );
  NOR2_X1 U117 ( .A1(n228), .A2(n229), .ZN(n225) );
  INV_X1 U118 ( .A(n200), .ZN(n229) );
  NAND4_X1 U119 ( .A1(n160), .A2(n152), .A3(n153), .A4(n141), .ZN(n144) );
  NAND2_X1 U120 ( .A1(n195), .A2(n197), .ZN(n211) );
  NAND4_X1 U121 ( .A1(n297), .A2(n51), .A3(n283), .A4(n56), .ZN(n189) );
  AOI21_X1 U122 ( .B1(n299), .B2(n298), .A(n300), .ZN(n297) );
  NOR2_X1 U123 ( .A1(n66), .A2(n304), .ZN(n302) );
  AOI21_X1 U124 ( .B1(n155), .B2(n153), .A(n156), .ZN(n150) );
  NAND2_X1 U125 ( .A1(n286), .A2(n8), .ZN(n325) );
  INV_X1 U126 ( .A(n289), .ZN(n287) );
  OAI21_X1 U127 ( .B1(n12), .B2(n342), .A(n337), .ZN(n341) );
  OAI21_X1 U128 ( .B1(n309), .B2(n310), .A(n278), .ZN(n308) );
  NAND2_X1 U129 ( .A1(n322), .A2(n277), .ZN(n321) );
  NAND2_X1 U130 ( .A1(n90), .A2(n85), .ZN(n295) );
  AND2_X1 U131 ( .A1(n171), .A2(n58), .ZN(n174) );
  AND2_X1 U132 ( .A1(n170), .A2(n159), .ZN(n58) );
  NAND2_X1 U133 ( .A1(n143), .A2(n140), .ZN(n116) );
  NOR2_X1 U134 ( .A1(n230), .A2(n231), .ZN(n228) );
  INV_X1 U135 ( .A(n206), .ZN(n230) );
  NAND2_X1 U136 ( .A1(n85), .A2(n86), .ZN(n84) );
  NAND2_X1 U137 ( .A1(n16), .A2(n88), .ZN(n86) );
  NAND2_X1 U138 ( .A1(n268), .A2(n263), .ZN(n267) );
  NAND2_X1 U139 ( .A1(n346), .A2(n72), .ZN(n343) );
  NAND2_X1 U140 ( .A1(n348), .A2(n349), .ZN(n346) );
  NOR2_X1 U141 ( .A1(n289), .A2(n296), .ZN(n290) );
  NAND2_X1 U142 ( .A1(n194), .A2(n195), .ZN(n113) );
  OAI21_X1 U143 ( .B1(n30), .B2(n61), .A(n196), .ZN(n194) );
  AND2_X1 U144 ( .A1(n197), .A2(n198), .ZN(n196) );
  NAND2_X1 U145 ( .A1(n157), .A2(n158), .ZN(n156) );
  NAND2_X1 U146 ( .A1(n204), .A2(n203), .ZN(n112) );
  NOR2_X1 U147 ( .A1(n187), .A2(n205), .ZN(n203) );
  NAND2_X1 U148 ( .A1(n330), .A2(n331), .ZN(n288) );
  AND2_X1 U149 ( .A1(n337), .A2(n338), .ZN(n330) );
  NAND2_X1 U150 ( .A1(n332), .A2(n333), .ZN(n331) );
  NAND2_X1 U151 ( .A1(n72), .A2(n335), .ZN(n332) );
  NAND2_X1 U152 ( .A1(n176), .A2(n9), .ZN(n171) );
  AND3_X1 U153 ( .A1(n120), .A2(n117), .A3(n118), .ZN(n59) );
  AND2_X1 U154 ( .A1(n279), .A2(n315), .ZN(n60) );
  NAND2_X1 U155 ( .A1(n274), .A2(n275), .ZN(n192) );
  AND2_X1 U156 ( .A1(n281), .A2(n282), .ZN(n274) );
  OAI211_X1 U157 ( .C1(n276), .C2(n277), .A(n278), .B(n279), .ZN(n275) );
  NAND2_X1 U158 ( .A1(n362), .A2(n363), .ZN(n293) );
  AND2_X1 U159 ( .A1(n94), .A2(n87), .ZN(n362) );
  INV_X1 U160 ( .A(A[0]), .ZN(n305) );
  NAND2_X1 U161 ( .A1(n173), .A2(n174), .ZN(n172) );
  AND2_X1 U162 ( .A1(n199), .A2(n200), .ZN(n61) );
  OAI21_X1 U163 ( .B1(n121), .B2(n122), .A(n123), .ZN(n119) );
  NAND2_X1 U164 ( .A1(n117), .A2(n118), .ZN(n115) );
  NAND2_X1 U165 ( .A1(n89), .A2(n90), .ZN(n83) );
  NAND2_X1 U166 ( .A1(n141), .A2(n157), .ZN(n164) );
  NAND2_X1 U167 ( .A1(n191), .A2(n38), .ZN(n307) );
  NAND2_X1 U168 ( .A1(n286), .A2(n338), .ZN(n340) );
  NAND2_X1 U169 ( .A1(n140), .A2(n138), .ZN(n147) );
  INV_X1 U170 ( .A(n199), .ZN(n217) );
  INV_X1 U171 ( .A(A[26]), .ZN(n178) );
  INV_X1 U172 ( .A(B[12]), .ZN(n339) );
  INV_X1 U173 ( .A(A[27]), .ZN(n166) );
  INV_X1 U174 ( .A(B[14]), .ZN(n313) );
  INV_X1 U175 ( .A(B[6]), .ZN(n360) );
  NAND2_X1 U176 ( .A1(A[21]), .A2(n223), .ZN(n199) );
  INV_X1 U177 ( .A(A[17]), .ZN(n240) );
  INV_X1 U178 ( .A(A[21]), .ZN(n224) );
  INV_X1 U179 ( .A(A[20]), .ZN(n247) );
  NAND2_X1 U180 ( .A1(A[20]), .A2(n246), .ZN(n200) );
  INV_X1 U181 ( .A(A[24]), .ZN(n209) );
  INV_X1 U182 ( .A(B[13]), .ZN(n326) );
  INV_X1 U183 ( .A(B[5]), .ZN(n365) );
  INV_X1 U184 ( .A(A[22]), .ZN(n221) );
  INV_X1 U185 ( .A(A[28]), .ZN(n162) );
  NAND2_X1 U186 ( .A1(B[7]), .A2(n359), .ZN(n89) );
  NAND2_X1 U187 ( .A1(B[25]), .A2(n183), .ZN(n152) );
  INV_X1 U188 ( .A(A[25]), .ZN(n183) );
  NAND2_X1 U189 ( .A1(B[6]), .A2(n367), .ZN(n87) );
  NAND2_X1 U190 ( .A1(A[26]), .A2(n177), .ZN(n158) );
  INV_X1 U191 ( .A(B[11]), .ZN(n344) );
  INV_X1 U192 ( .A(A[23]), .ZN(n213) );
  NAND2_X1 U193 ( .A1(A[27]), .A2(n165), .ZN(n157) );
  NAND2_X1 U194 ( .A1(A[18]), .A2(n264), .ZN(n242) );
  NAND2_X1 U195 ( .A1(B[14]), .A2(n314), .ZN(n282) );
  NAND2_X1 U196 ( .A1(B[5]), .A2(n366), .ZN(n94) );
  NAND2_X1 U197 ( .A1(A[22]), .A2(n220), .ZN(n198) );
  INV_X1 U198 ( .A(A[19]), .ZN(n255) );
  INV_X1 U199 ( .A(A[18]), .ZN(n265) );
  NAND2_X1 U200 ( .A1(A[23]), .A2(n212), .ZN(n197) );
  NAND2_X1 U201 ( .A1(A[28]), .A2(n161), .ZN(n138) );
  NAND2_X1 U202 ( .A1(B[17]), .A2(n240), .ZN(n244) );
  NAND2_X1 U203 ( .A1(A[19]), .A2(n254), .ZN(n243) );
  INV_X1 U204 ( .A(B[10]), .ZN(n370) );
  INV_X1 U205 ( .A(B[7]), .ZN(n361) );
  NOR2_X1 U206 ( .A1(B[17]), .A2(n240), .ZN(n238) );
  INV_X1 U207 ( .A(A[16]), .ZN(n241) );
  NAND2_X1 U208 ( .A1(n258), .A2(n257), .ZN(n253) );
  NOR2_X1 U209 ( .A1(n260), .A2(n261), .ZN(n257) );
  INV_X1 U210 ( .A(n262), .ZN(n261) );
  INV_X1 U211 ( .A(B[8]), .ZN(n336) );
  NAND2_X1 U212 ( .A1(A[25]), .A2(n182), .ZN(n159) );
  INV_X1 U213 ( .A(B[25]), .ZN(n182) );
  NAND2_X1 U214 ( .A1(n235), .A2(n236), .ZN(n204) );
  AND2_X1 U215 ( .A1(n242), .A2(n243), .ZN(n235) );
  NAND2_X1 U216 ( .A1(B[8]), .A2(n368), .ZN(n74) );
  INV_X1 U217 ( .A(A[29]), .ZN(n146) );
  INV_X1 U218 ( .A(A[30]), .ZN(n129) );
  NAND2_X1 U219 ( .A1(A[16]), .A2(n271), .ZN(n263) );
  NAND2_X1 U220 ( .A1(A[17]), .A2(n259), .ZN(n262) );
  NAND2_X1 U221 ( .A1(A[29]), .A2(n145), .ZN(n122) );
  AOI21_X1 U222 ( .B1(B[17]), .B2(n240), .A(n263), .ZN(n260) );
  NAND2_X1 U223 ( .A1(B[17]), .A2(n240), .ZN(n269) );
  NAND2_X1 U224 ( .A1(A[30]), .A2(n130), .ZN(n123) );
  INV_X1 U225 ( .A(B[17]), .ZN(n259) );
  XOR2_X1 U226 ( .A(B[31]), .B(A[31]), .Z(n62) );
  NAND2_X1 U227 ( .A1(n138), .A2(n139), .ZN(n120) );
  NAND2_X1 U228 ( .A1(A[0]), .A2(n65), .ZN(n249) );
  NAND2_X1 U229 ( .A1(n190), .A2(n188), .ZN(n285) );
  NAND2_X1 U230 ( .A1(n204), .A2(n207), .ZN(n231) );
  NAND2_X1 U231 ( .A1(n207), .A2(n243), .ZN(n250) );
  NOR2_X1 U232 ( .A1(n285), .A2(n27), .ZN(n272) );
  NAND2_X1 U233 ( .A1(B[4]), .A2(n358), .ZN(n99) );
  INV_X1 U234 ( .A(B[4]), .ZN(n364) );
  NAND2_X1 U235 ( .A1(n334), .A2(n337), .ZN(n345) );
  NAND2_X1 U236 ( .A1(B[10]), .A2(n371), .ZN(n334) );
  NAND2_X1 U237 ( .A1(n354), .A2(n105), .ZN(n298) );
  XNOR2_X1 U238 ( .A(n42), .B(n270), .ZN(DIFF[16]) );
  NAND2_X1 U239 ( .A1(n226), .A2(n42), .ZN(n234) );
  NAND2_X1 U240 ( .A1(n15), .A2(n72), .ZN(n70) );
  AND2_X1 U241 ( .A1(n71), .A2(n334), .ZN(n333) );
  AND2_X1 U242 ( .A1(n71), .A2(n74), .ZN(n348) );
  INV_X1 U243 ( .A(B[29]), .ZN(n145) );
  NAND2_X1 U244 ( .A1(B[29]), .A2(n146), .ZN(n118) );
  INV_X1 U245 ( .A(B[23]), .ZN(n212) );
  NAND2_X1 U246 ( .A1(B[23]), .A2(n213), .ZN(n195) );
  NAND2_X1 U247 ( .A1(n150), .A2(n151), .ZN(n142) );
  NAND2_X1 U248 ( .A1(B[19]), .A2(n255), .ZN(n207) );
  INV_X1 U249 ( .A(B[19]), .ZN(n254) );
  OAI21_X1 U250 ( .B1(n185), .B2(n186), .A(n43), .ZN(n114) );
  NAND2_X1 U251 ( .A1(B[26]), .A2(n178), .ZN(n153) );
  INV_X1 U252 ( .A(B[26]), .ZN(n177) );
  NAND2_X1 U253 ( .A1(n48), .A2(n365), .ZN(n93) );
  INV_X1 U254 ( .A(A[5]), .ZN(n366) );
  NAND2_X1 U255 ( .A1(n108), .A2(n109), .ZN(n107) );
  INV_X1 U256 ( .A(A[3]), .ZN(n357) );
  NAND2_X1 U257 ( .A1(A[3]), .A2(n356), .ZN(n106) );
  NAND2_X1 U258 ( .A1(n29), .A2(n99), .ZN(n100) );
  NAND2_X1 U259 ( .A1(n93), .A2(n98), .ZN(n363) );
  NAND2_X1 U260 ( .A1(A[11]), .A2(n344), .ZN(n338) );
  XNOR2_X1 U261 ( .A(n184), .B(n19), .ZN(DIFF[24]) );
  NAND2_X1 U262 ( .A1(A[12]), .A2(n339), .ZN(n277) );
  NAND2_X1 U263 ( .A1(A[15]), .A2(n312), .ZN(n191) );
  INV_X1 U264 ( .A(A[15]), .ZN(n311) );
  NAND2_X1 U265 ( .A1(B[27]), .A2(n166), .ZN(n141) );
  INV_X1 U266 ( .A(B[27]), .ZN(n165) );
  NAND2_X1 U267 ( .A1(A[4]), .A2(n364), .ZN(n98) );
  INV_X1 U268 ( .A(A[4]), .ZN(n358) );
  NAND4_X1 U269 ( .A1(n206), .A2(n201), .A3(n202), .A4(n195), .ZN(n187) );
  NAND2_X1 U270 ( .A1(n217), .A2(n202), .ZN(n214) );
  NAND2_X1 U271 ( .A1(n202), .A2(n198), .ZN(n219) );
  INV_X1 U272 ( .A(n227), .ZN(n226) );
  NAND2_X1 U273 ( .A1(A[9]), .A2(n347), .ZN(n72) );
  OAI211_X1 U274 ( .C1(n237), .C2(n238), .A(n244), .B(n239), .ZN(n236) );
  NAND2_X1 U275 ( .A1(n239), .A2(n242), .ZN(n256) );
  INV_X1 U276 ( .A(A[1]), .ZN(n304) );
  NAND2_X1 U277 ( .A1(n1), .A2(n360), .ZN(n85) );
  INV_X1 U278 ( .A(A[6]), .ZN(n367) );
  NAND2_X1 U279 ( .A1(A[14]), .A2(n313), .ZN(n278) );
  INV_X1 U280 ( .A(A[14]), .ZN(n314) );
  NAND2_X1 U281 ( .A1(A[13]), .A2(n326), .ZN(n279) );
  INV_X1 U282 ( .A(A[13]), .ZN(n327) );
  NAND2_X1 U283 ( .A1(A[7]), .A2(n361), .ZN(n90) );
  INV_X1 U284 ( .A(A[7]), .ZN(n359) );
  INV_X1 U285 ( .A(B[20]), .ZN(n246) );
  NAND2_X1 U286 ( .A1(B[20]), .A2(n247), .ZN(n206) );
  NAND4_X1 U287 ( .A1(n244), .A2(n245), .A3(n239), .A4(n207), .ZN(n227) );
  NAND2_X1 U288 ( .A1(n245), .A2(n42), .ZN(n268) );
  NAND2_X1 U289 ( .A1(n263), .A2(n245), .ZN(n270) );
  INV_X1 U290 ( .A(B[28]), .ZN(n161) );
  NAND2_X1 U291 ( .A1(B[28]), .A2(n162), .ZN(n140) );
  INV_X1 U292 ( .A(B[21]), .ZN(n223) );
  NAND2_X1 U293 ( .A1(B[21]), .A2(n224), .ZN(n201) );
  INV_X1 U294 ( .A(B[15]), .ZN(n312) );
  NAND2_X1 U295 ( .A1(B[15]), .A2(n311), .ZN(n281) );
  INV_X1 U296 ( .A(B[22]), .ZN(n220) );
  NAND2_X1 U297 ( .A1(B[22]), .A2(n221), .ZN(n202) );
  INV_X1 U298 ( .A(B[18]), .ZN(n264) );
  NAND2_X1 U299 ( .A1(B[18]), .A2(n265), .ZN(n239) );
  INV_X1 U300 ( .A(B[9]), .ZN(n347) );
  NAND2_X1 U301 ( .A1(B[24]), .A2(n209), .ZN(n160) );
  NAND2_X1 U302 ( .A1(n6), .A2(n370), .ZN(n337) );
  INV_X1 U303 ( .A(A[10]), .ZN(n371) );
  INV_X1 U304 ( .A(B[30]), .ZN(n130) );
  NAND2_X1 U305 ( .A1(B[30]), .A2(n129), .ZN(n117) );
  NAND2_X1 U306 ( .A1(n160), .A2(n154), .ZN(n184) );
  NAND2_X1 U307 ( .A1(n112), .A2(n154), .ZN(n176) );
  NAND2_X1 U308 ( .A1(A[8]), .A2(n336), .ZN(n335) );
  INV_X1 U309 ( .A(A[8]), .ZN(n368) );
  NAND2_X1 U310 ( .A1(B[9]), .A2(n369), .ZN(n71) );
  INV_X1 U311 ( .A(A[9]), .ZN(n369) );
  AND2_X1 U312 ( .A1(n50), .A2(n355), .ZN(n63) );
  INV_X1 U313 ( .A(A[2]), .ZN(n355) );
  NAND2_X1 U314 ( .A1(n66), .A2(n304), .ZN(n303) );
  OAI21_X1 U315 ( .B1(n33), .B2(n181), .A(n154), .ZN(n180) );
  OAI21_X1 U316 ( .B1(n33), .B2(n144), .A(n149), .ZN(n148) );
  OAI21_X1 U317 ( .B1(n33), .B2(n116), .A(n137), .ZN(n136) );
  OAI21_X1 U318 ( .B1(n33), .B2(n125), .A(n126), .ZN(n124) );
  NAND2_X1 U319 ( .A1(n249), .A2(n351), .ZN(DIFF[0]) );
  INV_X1 U320 ( .A(B[16]), .ZN(n271) );
  NAND2_X1 U321 ( .A1(B[16]), .A2(n241), .ZN(n245) );
  NOR2_X1 U322 ( .A1(B[16]), .A2(n241), .ZN(n237) );
  NAND2_X1 U323 ( .A1(n303), .A2(n133), .ZN(n248) );
  NAND2_X1 U324 ( .A1(n64), .A2(n305), .ZN(n351) );
  NOR2_X1 U325 ( .A1(n64), .A2(n305), .ZN(n301) );
  NAND2_X1 U326 ( .A1(n135), .A2(n103), .ZN(n131) );
  NAND2_X1 U327 ( .A1(A[2]), .A2(n68), .ZN(n103) );
  OAI211_X1 U328 ( .C1(n301), .C2(n302), .A(n303), .B(n135), .ZN(n299) );
  OAI21_X1 U329 ( .B1(n50), .B2(n355), .A(n106), .ZN(n354) );
  NAND2_X1 U330 ( .A1(n50), .A2(n355), .ZN(n135) );
  OAI211_X1 U331 ( .C1(A[17]), .C2(n259), .A(n25), .B(n245), .ZN(n258) );
  XNOR2_X1 U332 ( .A(n210), .B(n211), .ZN(DIFF[23]) );
  OAI21_X1 U333 ( .B1(n132), .B2(n55), .A(n133), .ZN(n104) );
  INV_X1 U334 ( .A(B[24]), .ZN(n208) );
  XNOR2_X1 U335 ( .A(n62), .B(n107), .ZN(DIFF[31]) );
  OAI21_X1 U336 ( .B1(n168), .B2(n44), .A(n153), .ZN(n167) );
  NAND2_X1 U337 ( .A1(n167), .A2(n32), .ZN(n163) );
  XNOR2_X1 U338 ( .A(n216), .B(n222), .ZN(DIFF[21]) );
  NAND2_X1 U339 ( .A1(n17), .A2(n225), .ZN(n216) );
  NAND2_X1 U340 ( .A1(n291), .A2(n290), .ZN(n190) );
  AOI21_X1 U341 ( .B1(n292), .B2(n293), .A(n294), .ZN(n291) );
  NAND2_X1 U342 ( .A1(A[1]), .A2(n67), .ZN(n133) );
  NAND2_X1 U343 ( .A1(B[3]), .A2(n357), .ZN(n105) );
  INV_X1 U344 ( .A(B[3]), .ZN(n356) );
  XNOR2_X1 U345 ( .A(n37), .B(n100), .ZN(DIFF[4]) );
  AOI21_X1 U346 ( .B1(n56), .B2(n37), .A(n82), .ZN(n78) );
  NAND2_X1 U347 ( .A1(n56), .A2(n81), .ZN(n77) );
  NAND2_X1 U348 ( .A1(n81), .A2(n99), .ZN(n97) );
  NAND2_X1 U349 ( .A1(n56), .A2(n37), .ZN(n324) );
  NAND4_X1 U350 ( .A1(n52), .A2(n51), .A3(n283), .A4(n56), .ZN(n193) );
  INV_X1 U351 ( .A(B[1]), .ZN(n67) );
  XNOR2_X1 U352 ( .A(n163), .B(n164), .ZN(DIFF[27]) );
  XNOR2_X1 U353 ( .A(n218), .B(n219), .ZN(DIFF[22]) );
  INV_X1 U354 ( .A(n65), .ZN(n64) );
  INV_X1 U355 ( .A(B[0]), .ZN(n65) );
  INV_X1 U356 ( .A(n67), .ZN(n66) );
  INV_X1 U357 ( .A(B[2]), .ZN(n68) );
  NOR2_X1 U358 ( .A1(n75), .A2(n80), .ZN(n79) );
  INV_X1 U359 ( .A(n74), .ZN(n80) );
  INV_X1 U360 ( .A(n335), .ZN(n75) );
  XNOR2_X1 U361 ( .A(n88), .B(n91), .ZN(DIFF[6]) );
  INV_X1 U362 ( .A(n94), .ZN(n92) );
  OAI21_X1 U363 ( .B1(n102), .B2(n63), .A(n103), .ZN(n101) );
  INV_X1 U364 ( .A(n104), .ZN(n102) );
  NAND3_X1 U365 ( .A1(n114), .A2(n113), .A3(n112), .ZN(n111) );
  INV_X1 U366 ( .A(n117), .ZN(n121) );
  INV_X1 U367 ( .A(n122), .ZN(n127) );
  NAND2_X1 U368 ( .A1(n118), .A2(n128), .ZN(n125) );
  INV_X1 U369 ( .A(n116), .ZN(n128) );
  XNOR2_X1 U370 ( .A(n131), .B(n104), .ZN(DIFF[2]) );
  INV_X1 U371 ( .A(n134), .ZN(n132) );
  INV_X1 U372 ( .A(n120), .ZN(n137) );
  NAND3_X1 U373 ( .A1(n142), .A2(n141), .A3(n140), .ZN(n139) );
  INV_X1 U374 ( .A(n144), .ZN(n143) );
  XNOR2_X1 U375 ( .A(n148), .B(n147), .ZN(DIFF[28]) );
  NAND3_X1 U376 ( .A1(n152), .A2(n36), .A3(n153), .ZN(n151) );
  INV_X1 U377 ( .A(n159), .ZN(n155) );
  NAND3_X1 U378 ( .A1(n171), .A2(n159), .A3(n170), .ZN(n168) );
  INV_X1 U379 ( .A(n113), .ZN(n175) );
  NAND3_X1 U380 ( .A1(n42), .A2(n9), .A3(n43), .ZN(n173) );
  XNOR2_X1 U381 ( .A(n179), .B(n180), .ZN(DIFF[25]) );
  INV_X1 U382 ( .A(n160), .ZN(n181) );
  NAND3_X1 U383 ( .A1(n188), .A2(n189), .A3(n190), .ZN(n186) );
  NAND3_X1 U384 ( .A1(n193), .A2(n192), .A3(n191), .ZN(n185) );
  INV_X1 U385 ( .A(n207), .ZN(n205) );
  NAND3_X1 U386 ( .A1(n215), .A2(n214), .A3(n198), .ZN(n210) );
  XNOR2_X1 U387 ( .A(n251), .B(n250), .ZN(DIFF[19]) );
  OAI21_X1 U388 ( .B1(n20), .B2(n252), .A(n242), .ZN(n251) );
  INV_X1 U389 ( .A(n239), .ZN(n252) );
  INV_X1 U390 ( .A(n280), .ZN(n276) );
  NAND3_X1 U391 ( .A1(n288), .A2(n287), .A3(n286), .ZN(n188) );
  INV_X1 U392 ( .A(n89), .ZN(n294) );
  INV_X1 U393 ( .A(n295), .ZN(n292) );
  INV_X1 U394 ( .A(n296), .ZN(n283) );
  XNOR2_X1 U395 ( .A(n308), .B(n307), .ZN(DIFF[15]) );
  INV_X1 U396 ( .A(n282), .ZN(n310) );
  INV_X1 U397 ( .A(n277), .ZN(n316) );
  NAND3_X1 U398 ( .A1(n318), .A2(n306), .A3(n319), .ZN(n322) );
  XNOR2_X1 U399 ( .A(n328), .B(n329), .ZN(DIFF[12]) );
  INV_X1 U400 ( .A(n76), .ZN(n82) );
  XNOR2_X1 U401 ( .A(n340), .B(n341), .ZN(DIFF[11]) );
  INV_X1 U402 ( .A(n334), .ZN(n342) );
  NAND3_X1 U403 ( .A1(n35), .A2(n105), .A3(n350), .ZN(n284) );
  NOR2_X1 U404 ( .A1(n300), .A2(n63), .ZN(n353) );
  INV_X1 U405 ( .A(n105), .ZN(n300) );
endmodule


module ALU_N32_DW01_cmp6_4 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  XNOR2_X1 U1 ( .A(B[17]), .B(A[17]), .ZN(n23) );
  XNOR2_X1 U2 ( .A(B[25]), .B(A[25]), .ZN(n13) );
  XNOR2_X1 U3 ( .A(B[0]), .B(A[0]), .ZN(n34) );
  XNOR2_X1 U4 ( .A(B[31]), .B(A[31]), .ZN(n7) );
  XNOR2_X1 U5 ( .A(B[29]), .B(A[29]), .ZN(n9) );
  XNOR2_X1 U6 ( .A(B[23]), .B(A[23]), .ZN(n17) );
  XNOR2_X1 U7 ( .A(B[26]), .B(A[26]), .ZN(n12) );
  XNOR2_X1 U8 ( .A(B[5]), .B(A[5]), .ZN(n29) );
  XNOR2_X1 U9 ( .A(B[11]), .B(A[11]), .ZN(n41) );
  XNOR2_X1 U10 ( .A(B[12]), .B(A[12]), .ZN(n40) );
  XNOR2_X1 U11 ( .A(B[27]), .B(A[27]), .ZN(n11) );
  XNOR2_X1 U12 ( .A(B[4]), .B(A[4]), .ZN(n30) );
  XNOR2_X1 U13 ( .A(B[19]), .B(A[19]), .ZN(n21) );
  XNOR2_X1 U14 ( .A(B[6]), .B(A[6]), .ZN(n28) );
  XNOR2_X1 U15 ( .A(B[14]), .B(A[14]), .ZN(n38) );
  XNOR2_X1 U16 ( .A(B[13]), .B(A[13]), .ZN(n39) );
  XNOR2_X1 U17 ( .A(B[7]), .B(A[7]), .ZN(n27) );
  XNOR2_X1 U18 ( .A(B[20]), .B(A[20]), .ZN(n20) );
  XNOR2_X1 U19 ( .A(B[28]), .B(A[28]), .ZN(n10) );
  XNOR2_X1 U20 ( .A(B[21]), .B(A[21]), .ZN(n19) );
  XNOR2_X1 U21 ( .A(B[15]), .B(A[15]), .ZN(n37) );
  XNOR2_X1 U22 ( .A(B[22]), .B(A[22]), .ZN(n18) );
  XNOR2_X1 U23 ( .A(B[18]), .B(A[18]), .ZN(n22) );
  XNOR2_X1 U24 ( .A(B[9]), .B(A[9]), .ZN(n43) );
  XNOR2_X1 U25 ( .A(B[24]), .B(A[24]), .ZN(n14) );
  XNOR2_X1 U26 ( .A(B[10]), .B(A[10]), .ZN(n42) );
  XNOR2_X1 U27 ( .A(B[30]), .B(A[30]), .ZN(n8) );
  XNOR2_X1 U28 ( .A(B[8]), .B(A[8]), .ZN(n44) );
  XNOR2_X1 U29 ( .A(B[16]), .B(A[16]), .ZN(n24) );
  XNOR2_X1 U30 ( .A(B[1]), .B(A[1]), .ZN(n32) );
  XNOR2_X1 U31 ( .A(B[2]), .B(A[2]), .ZN(n33) );
  XNOR2_X1 U32 ( .A(B[3]), .B(A[3]), .ZN(n31) );
  NAND4_X1 U33 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(NE) );
  NOR2_X1 U34 ( .A1(n5), .A2(n6), .ZN(n4) );
  NAND4_X1 U35 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n6) );
  NAND4_X1 U36 ( .A1(n11), .A2(n12), .A3(n13), .A4(n14), .ZN(n5) );
  NOR2_X1 U37 ( .A1(n15), .A2(n16), .ZN(n3) );
  NAND4_X1 U38 ( .A1(n17), .A2(n18), .A3(n19), .A4(n20), .ZN(n16) );
  NAND4_X1 U39 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n15) );
  NOR2_X1 U40 ( .A1(n25), .A2(n26), .ZN(n2) );
  NAND4_X1 U41 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(n26) );
  NAND4_X1 U42 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(n25) );
  NOR2_X1 U43 ( .A1(n35), .A2(n36), .ZN(n1) );
  NAND4_X1 U44 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n36) );
  NAND4_X1 U45 ( .A1(n41), .A2(n42), .A3(n43), .A4(n44), .ZN(n35) );
endmodule


module ALU_N32_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   net46653, net46652, net46632, net46631, net46630, net46626, net46601,
         net46600, net46590, net46588, net46579, net46575, net46571, net46570,
         net46569, net46568, net46564, net46562, net46561, net46556, net46553,
         net46546, net46536, net46535, net46527, net46523, net46522, net46506,
         net46496, net46490, net46488, net46481, net46480, net46479, net46478,
         net46469, net46467, net46456, net46455, net46454, net46452, net46451,
         net46450, net46444, net46443, net46442, net46439, net46436, net46413,
         net46412, net46404, net46360, net46358, net46355, net46354, net46352,
         net46346, net46307, net46304, net46303, net46301, net46277, net52114,
         net52555, net52600, net52631, net52658, net52679, net52700, net52718,
         net52836, net52904, net52925, net52944, net46560, net46559, net46555,
         net46552, net46549, net46357, net46529, net46462, net46460, net46459,
         net46453, net46438, net52107, net46550, net46548, net46486, net46484,
         net46475, net46406, net46362, net46353, net46321, net46278, net52652,
         net52544, net52111, net46563, net46558, net46557, net46551, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242;

  OR2_X1 U2 ( .A1(B[3]), .A2(A[3]), .ZN(net46303) );
  INV_X1 U3 ( .A(net52925), .ZN(n1) );
  CLKBUF_X1 U4 ( .A(A[7]), .Z(n2) );
  OR2_X2 U5 ( .A1(B[25]), .A2(A[25]), .ZN(n134) );
  AND2_X1 U6 ( .A1(A[6]), .A2(B[6]), .ZN(n38) );
  BUF_X1 U7 ( .A(net52544), .Z(n3) );
  CLKBUF_X1 U8 ( .A(A[9]), .Z(n4) );
  CLKBUF_X1 U9 ( .A(A[7]), .Z(n5) );
  AND3_X1 U10 ( .A1(net46535), .A2(net46536), .A3(net46626), .ZN(n6) );
  AND2_X1 U11 ( .A1(net46354), .A2(net46355), .ZN(n7) );
  OR2_X1 U12 ( .A1(n91), .A2(n90), .ZN(n8) );
  OR2_X1 U13 ( .A1(n91), .A2(n101), .ZN(n9) );
  INV_X1 U14 ( .A(n40), .ZN(n73) );
  OR2_X1 U15 ( .A1(B[24]), .A2(A[24]), .ZN(n142) );
  CLKBUF_X1 U16 ( .A(B[9]), .Z(n10) );
  CLKBUF_X1 U17 ( .A(net46601), .Z(n11) );
  AND2_X1 U18 ( .A1(net46630), .A2(n38), .ZN(n12) );
  INV_X1 U19 ( .A(n38), .ZN(n67) );
  CLKBUF_X1 U20 ( .A(B[22]), .Z(n13) );
  CLKBUF_X1 U21 ( .A(A[12]), .Z(n14) );
  CLKBUF_X1 U22 ( .A(net46563), .Z(n15) );
  OR2_X2 U23 ( .A1(B[14]), .A2(A[14]), .ZN(net46553) );
  CLKBUF_X1 U24 ( .A(n228), .Z(n16) );
  CLKBUF_X1 U25 ( .A(B[7]), .Z(n17) );
  BUF_X1 U26 ( .A(B[3]), .Z(n47) );
  OR2_X1 U27 ( .A1(B[27]), .A2(A[27]), .ZN(n127) );
  INV_X1 U28 ( .A(n78), .ZN(n18) );
  OR2_X1 U29 ( .A1(A[2]), .A2(B[2]), .ZN(n108) );
  INV_X1 U30 ( .A(net52631), .ZN(net46523) );
  OR2_X1 U31 ( .A1(A[12]), .A2(B[12]), .ZN(net46563) );
  NOR2_X1 U32 ( .A1(n17), .A2(n5), .ZN(n19) );
  AND3_X1 U33 ( .A1(net46562), .A2(net46561), .A3(net52700), .ZN(net52944) );
  NAND4_X1 U34 ( .A1(n27), .A2(net52700), .A3(n31), .A4(net52904), .ZN(n20) );
  AND2_X1 U35 ( .A1(n127), .A2(n134), .ZN(n21) );
  OR2_X1 U36 ( .A1(B[18]), .A2(A[18]), .ZN(net46480) );
  AND2_X1 U37 ( .A1(net46481), .A2(net46480), .ZN(n178) );
  AND2_X1 U38 ( .A1(net52111), .A2(net52544), .ZN(net52652) );
  AOI21_X1 U39 ( .B1(net52652), .B2(net46486), .A(net46362), .ZN(net46484) );
  AND4_X1 U40 ( .A1(net46563), .A2(net46551), .A3(net46553), .A4(net46552), 
        .ZN(net52111) );
  AND2_X1 U41 ( .A1(net46600), .A2(net46601), .ZN(net52544) );
  NAND2_X1 U42 ( .A1(net52700), .A2(net52904), .ZN(net46490) );
  OR2_X1 U43 ( .A1(B[15]), .A2(A[15]), .ZN(net46551) );
  AND4_X1 U44 ( .A1(net46551), .A2(net46563), .A3(net46564), .A4(net46553), 
        .ZN(net52700) );
  INV_X1 U45 ( .A(net46551), .ZN(net46550) );
  CLKBUF_X1 U46 ( .A(net46551), .Z(net52555) );
  NAND2_X1 U47 ( .A1(net46557), .A2(net46558), .ZN(net46564) );
  INV_X1 U48 ( .A(A[13]), .ZN(net46558) );
  NAND2_X1 U49 ( .A1(net46557), .A2(net46558), .ZN(net46552) );
  INV_X1 U50 ( .A(B[13]), .ZN(net46557) );
  NAND2_X1 U51 ( .A1(n15), .A2(net46579), .ZN(net46590) );
  INV_X1 U52 ( .A(net46563), .ZN(net46588) );
  AND2_X1 U53 ( .A1(net46600), .A2(net46601), .ZN(net52904) );
  CLKBUF_X1 U54 ( .A(net46600), .Z(net52718) );
  NAND2_X1 U55 ( .A1(B[15]), .A2(A[15]), .ZN(net46559) );
  NAND2_X1 U56 ( .A1(B[13]), .A2(A[13]), .ZN(net46556) );
  NAND2_X1 U57 ( .A1(B[14]), .A2(A[14]), .ZN(net46560) );
  NAND2_X1 U58 ( .A1(B[12]), .A2(n14), .ZN(net46579) );
  NAND2_X1 U59 ( .A1(A[12]), .A2(B[12]), .ZN(net46555) );
  NOR2_X1 U60 ( .A1(net46321), .A2(net46353), .ZN(n22) );
  OAI21_X1 U61 ( .B1(n22), .B2(net46453), .A(net46462), .ZN(net46460) );
  INV_X1 U62 ( .A(net46406), .ZN(net46321) );
  OAI21_X1 U63 ( .B1(net46475), .B2(net52944), .A(net52107), .ZN(net46406) );
  NAND2_X1 U64 ( .A1(net46354), .A2(net46355), .ZN(net46353) );
  NOR2_X1 U65 ( .A1(net46353), .A2(n1), .ZN(net46307) );
  AOI21_X1 U66 ( .B1(net52107), .B2(net46352), .A(net46353), .ZN(net46346) );
  NAND2_X1 U67 ( .A1(net46484), .A2(net46357), .ZN(net46475) );
  OAI21_X1 U68 ( .B1(net46475), .B2(net52944), .A(net52107), .ZN(net52925) );
  AOI21_X1 U69 ( .B1(net46548), .B2(net46549), .A(net46550), .ZN(net46362) );
  AOI21_X1 U70 ( .B1(net46549), .B2(net46548), .A(net46550), .ZN(net52658) );
  AND2_X1 U71 ( .A1(net46559), .A2(net46560), .ZN(net46548) );
  NAND2_X1 U72 ( .A1(n23), .A2(net46488), .ZN(net46486) );
  NOR2_X1 U73 ( .A1(net52600), .A2(net46278), .ZN(n23) );
  INV_X1 U74 ( .A(net46536), .ZN(net46278) );
  NOR2_X1 U75 ( .A1(n12), .A2(net46278), .ZN(net46529) );
  NOR2_X1 U76 ( .A1(net46278), .A2(n19), .ZN(net46277) );
  AND4_X1 U77 ( .A1(net46478), .A2(net46479), .A3(net46480), .A4(net46481), 
        .ZN(net52107) );
  AOI21_X1 U78 ( .B1(net46354), .B2(net46355), .A(net46412), .ZN(net46413) );
  INV_X1 U79 ( .A(net46355), .ZN(net46506) );
  AND3_X2 U80 ( .A1(net46527), .A2(n20), .A3(net46358), .ZN(net52631) );
  XNOR2_X1 U81 ( .A(net46460), .B(net46459), .ZN(SUM[22]) );
  NAND2_X1 U82 ( .A1(net46444), .A2(net46438), .ZN(net46459) );
  NOR2_X1 U83 ( .A1(n25), .A2(n26), .ZN(net46462) );
  NOR2_X1 U84 ( .A1(net46453), .A2(net46442), .ZN(n26) );
  INV_X1 U85 ( .A(n24), .ZN(n25) );
  OR2_X1 U86 ( .A1(B[22]), .A2(A[22]), .ZN(net46444) );
  NAND2_X1 U87 ( .A1(B[22]), .A2(A[22]), .ZN(net46438) );
  INV_X1 U88 ( .A(net46438), .ZN(net46436) );
  OAI21_X1 U89 ( .B1(net46452), .B2(n24), .A(net46438), .ZN(net46451) );
  NAND2_X1 U90 ( .A1(net46443), .A2(net46439), .ZN(net46453) );
  NOR2_X1 U91 ( .A1(net46453), .A2(net46454), .ZN(net46450) );
  INV_X1 U92 ( .A(net46453), .ZN(net46456) );
  NAND2_X1 U93 ( .A1(B[20]), .A2(A[20]), .ZN(net46442) );
  NAND2_X1 U94 ( .A1(B[21]), .A2(A[21]), .ZN(n24) );
  NAND2_X1 U95 ( .A1(net46439), .A2(n24), .ZN(net46467) );
  AND2_X1 U96 ( .A1(n24), .A2(net46442), .ZN(net52114) );
  CLKBUF_X1 U97 ( .A(net46559), .Z(net52679) );
  OAI21_X1 U98 ( .B1(net46569), .B2(net46570), .A(net46560), .ZN(net46568) );
  NAND2_X1 U99 ( .A1(net46560), .A2(net46553), .ZN(net46575) );
  AOI21_X1 U100 ( .B1(net46488), .B2(net46529), .A(net46490), .ZN(net46360) );
  NAND4_X1 U101 ( .A1(n27), .A2(n31), .A3(net52700), .A4(net52904), .ZN(
        net46357) );
  AND2_X1 U102 ( .A1(net46631), .A2(net46632), .ZN(n31) );
  NAND3_X1 U103 ( .A1(n33), .A2(net46546), .A3(n32), .ZN(n27) );
  AND2_X1 U104 ( .A1(n28), .A2(net46304), .ZN(n32) );
  NAND2_X1 U105 ( .A1(net46303), .A2(n30), .ZN(n28) );
  INV_X1 U106 ( .A(net46301), .ZN(n30) );
  NAND2_X1 U107 ( .A1(net46652), .A2(net46653), .ZN(n33) );
  NAND3_X1 U108 ( .A1(net46564), .A2(net46553), .A3(n29), .ZN(net46549) );
  NAND2_X1 U109 ( .A1(net46555), .A2(net46556), .ZN(n29) );
  AND2_X2 U110 ( .A1(n34), .A2(n35), .ZN(n152) );
  OR2_X1 U111 ( .A1(net52114), .A2(n140), .ZN(n34) );
  AND2_X1 U112 ( .A1(n136), .A2(n139), .ZN(n35) );
  OR2_X1 U113 ( .A1(B[8]), .A2(A[8]), .ZN(n58) );
  BUF_X1 U114 ( .A(A[3]), .Z(n46) );
  AND3_X2 U115 ( .A1(n202), .A2(n237), .A3(net46304), .ZN(n40) );
  INV_X1 U116 ( .A(n108), .ZN(n36) );
  OAI21_X1 U117 ( .B1(net52631), .B2(n190), .A(n191), .ZN(n37) );
  CLKBUF_X1 U118 ( .A(net46303), .Z(net52836) );
  NAND2_X1 U119 ( .A1(B[5]), .A2(n48), .ZN(n39) );
  OR2_X1 U120 ( .A1(B[1]), .A2(A[1]), .ZN(n106) );
  AND3_X1 U121 ( .A1(n21), .A2(n126), .A3(n142), .ZN(n41) );
  OR2_X1 U122 ( .A1(net46346), .A2(n111), .ZN(n42) );
  NAND2_X1 U123 ( .A1(n42), .A2(n112), .ZN(n110) );
  BUF_X1 U124 ( .A(A[5]), .Z(n48) );
  AND2_X1 U125 ( .A1(n71), .A2(n74), .ZN(net46631) );
  BUF_X1 U126 ( .A(B[0]), .Z(n43) );
  INV_X1 U127 ( .A(n43), .ZN(n44) );
  INV_X1 U128 ( .A(n132), .ZN(n45) );
  AND2_X1 U129 ( .A1(n38), .A2(net46630), .ZN(net52600) );
  OR2_X1 U130 ( .A1(A[5]), .A2(B[5]), .ZN(n71) );
  NAND3_X1 U131 ( .A1(n142), .A2(n126), .A3(n21), .ZN(n135) );
  INV_X1 U132 ( .A(n49), .ZN(n176) );
  AND2_X2 U133 ( .A1(n7), .A2(net52925), .ZN(n49) );
  XOR2_X1 U134 ( .A(net46575), .B(n50), .Z(SUM[14]) );
  AND2_X1 U135 ( .A1(n204), .A2(net46556), .ZN(n50) );
  AND2_X1 U136 ( .A1(n184), .A2(n239), .ZN(SUM[0]) );
  OR2_X1 U137 ( .A1(B[10]), .A2(A[10]), .ZN(n218) );
  NAND2_X1 U138 ( .A1(n141), .A2(n41), .ZN(n91) );
  AOI21_X1 U139 ( .B1(n84), .B2(n92), .A(n96), .ZN(n95) );
  AOI21_X1 U140 ( .B1(net46413), .B2(n148), .A(n154), .ZN(n145) );
  NOR2_X1 U141 ( .A1(n149), .A2(n150), .ZN(n146) );
  OAI21_X1 U142 ( .B1(net46307), .B2(n8), .A(n82), .ZN(n81) );
  AOI21_X1 U143 ( .B1(n84), .B2(n83), .A(n85), .ZN(n82) );
  INV_X1 U144 ( .A(net46360), .ZN(net46358) );
  NOR2_X1 U145 ( .A1(net52944), .A2(net52658), .ZN(n115) );
  NOR2_X1 U146 ( .A1(net52944), .A2(net52658), .ZN(net46527) );
  NAND2_X1 U147 ( .A1(n104), .A2(n105), .ZN(n79) );
  NAND2_X1 U148 ( .A1(n106), .A2(n107), .ZN(n104) );
  INV_X1 U149 ( .A(n184), .ZN(n107) );
  NAND2_X1 U150 ( .A1(n106), .A2(n105), .ZN(n183) );
  OAI21_X1 U151 ( .B1(n63), .B2(n64), .A(n65), .ZN(n61) );
  NAND2_X1 U152 ( .A1(n155), .A2(n142), .ZN(n168) );
  NAND2_X1 U153 ( .A1(n126), .A2(n130), .ZN(n156) );
  OAI21_X1 U154 ( .B1(n166), .B2(n152), .A(n155), .ZN(n160) );
  OAI21_X1 U155 ( .B1(n208), .B2(n209), .A(n210), .ZN(n205) );
  NAND2_X1 U156 ( .A1(n211), .A2(n6), .ZN(n209) );
  OAI21_X1 U157 ( .B1(net52631), .B2(n190), .A(n191), .ZN(n187) );
  NAND2_X1 U158 ( .A1(net46479), .A2(net46478), .ZN(n190) );
  AOI21_X1 U159 ( .B1(n192), .B2(net46479), .A(n193), .ZN(n191) );
  OAI21_X1 U160 ( .B1(n230), .B2(n231), .A(n55), .ZN(n228) );
  NAND2_X1 U161 ( .A1(n120), .A2(n119), .ZN(n84) );
  NOR2_X1 U162 ( .A1(n122), .A2(n121), .ZN(n120) );
  AOI21_X1 U163 ( .B1(n137), .B2(n41), .A(n138), .ZN(n119) );
  AND2_X1 U164 ( .A1(net46546), .A2(n28), .ZN(n237) );
  NAND2_X1 U165 ( .A1(net52555), .A2(net52679), .ZN(n203) );
  NAND2_X1 U166 ( .A1(net46564), .A2(net46553), .ZN(net46570) );
  NAND2_X1 U167 ( .A1(n45), .A2(n131), .ZN(n163) );
  NAND2_X1 U168 ( .A1(net46480), .A2(n182), .ZN(n189) );
  NAND2_X1 U169 ( .A1(net46552), .A2(net46556), .ZN(n206) );
  NAND2_X1 U170 ( .A1(n220), .A2(n218), .ZN(n229) );
  NAND2_X1 U171 ( .A1(net46479), .A2(n181), .ZN(n195) );
  OAI21_X1 U172 ( .B1(net52631), .B2(net46522), .A(n194), .ZN(n196) );
  NAND2_X1 U173 ( .A1(n54), .A2(n55), .ZN(n53) );
  NOR2_X1 U174 ( .A1(net52114), .A2(n140), .ZN(n137) );
  OAI21_X1 U175 ( .B1(n86), .B2(n87), .A(n88), .ZN(n85) );
  AOI21_X1 U176 ( .B1(n160), .B2(n45), .A(n161), .ZN(n159) );
  NAND4_X1 U177 ( .A1(net46439), .A2(net46443), .A3(n170), .A4(net46444), .ZN(
        n167) );
  NOR2_X1 U178 ( .A1(net46412), .A2(n155), .ZN(n154) );
  AOI21_X1 U179 ( .B1(n84), .B2(n102), .A(n113), .ZN(n112) );
  NAND2_X1 U180 ( .A1(net46561), .A2(net46562), .ZN(n211) );
  NAND2_X1 U181 ( .A1(n134), .A2(n126), .ZN(net46412) );
  NOR2_X1 U182 ( .A1(n152), .A2(n153), .ZN(n149) );
  NAND2_X1 U183 ( .A1(net46404), .A2(n142), .ZN(n153) );
  NOR2_X1 U184 ( .A1(net46571), .A2(n207), .ZN(net46569) );
  XNOR2_X1 U185 ( .A(net46590), .B(n212), .ZN(SUM[12]) );
  NAND2_X1 U186 ( .A1(n213), .A2(n211), .ZN(n212) );
  NAND2_X1 U187 ( .A1(n207), .A2(net46552), .ZN(n204) );
  XNOR2_X1 U188 ( .A(n59), .B(net46277), .ZN(SUM[7]) );
  AOI21_X1 U189 ( .B1(n60), .B2(n61), .A(n38), .ZN(n59) );
  XNOR2_X1 U190 ( .A(n62), .B(n61), .ZN(SUM[6]) );
  NAND2_X1 U191 ( .A1(n60), .A2(n67), .ZN(n62) );
  NAND2_X1 U192 ( .A1(net46631), .A2(net46632), .ZN(n200) );
  NAND2_X1 U193 ( .A1(n136), .A2(n170), .ZN(n171) );
  NAND2_X1 U194 ( .A1(n65), .A2(n70), .ZN(n234) );
  NAND2_X1 U195 ( .A1(net46436), .A2(n170), .ZN(n139) );
  NAND2_X1 U196 ( .A1(n98), .A2(n102), .ZN(n101) );
  NAND2_X1 U197 ( .A1(n97), .A2(n98), .ZN(n87) );
  NAND2_X1 U198 ( .A1(n99), .A2(n100), .ZN(n97) );
  NAND2_X1 U199 ( .A1(n92), .A2(n89), .ZN(n90) );
  NAND2_X1 U200 ( .A1(n141), .A2(n142), .ZN(n162) );
  NAND2_X1 U201 ( .A1(n38), .A2(net46630), .ZN(net46535) );
  NAND2_X1 U202 ( .A1(net46561), .A2(n219), .ZN(n226) );
  OAI21_X1 U203 ( .B1(n131), .B2(n151), .A(n130), .ZN(n150) );
  INV_X1 U204 ( .A(n126), .ZN(n151) );
  NAND2_X1 U205 ( .A1(n194), .A2(net46478), .ZN(n197) );
  NAND2_X1 U206 ( .A1(n65), .A2(n71), .ZN(n68) );
  XNOR2_X1 U207 ( .A(n56), .B(n57), .ZN(SUM[8]) );
  NAND2_X1 U208 ( .A1(n215), .A2(n58), .ZN(n56) );
  NAND2_X1 U209 ( .A1(B[1]), .A2(A[1]), .ZN(n105) );
  NOR2_X1 U210 ( .A1(net46506), .A2(net46496), .ZN(n186) );
  NAND2_X1 U211 ( .A1(n127), .A2(n125), .ZN(n144) );
  NAND2_X1 U212 ( .A1(n43), .A2(A[0]), .ZN(n184) );
  NAND2_X1 U213 ( .A1(n18), .A2(net46301), .ZN(n103) );
  NOR2_X1 U214 ( .A1(net46450), .A2(net46451), .ZN(n174) );
  NAND2_X1 U215 ( .A1(n98), .A2(n100), .ZN(n109) );
  NAND2_X1 U216 ( .A1(net52836), .A2(net46304), .ZN(n75) );
  NAND2_X1 U217 ( .A1(n99), .A2(n102), .ZN(n116) );
  NAND2_X1 U218 ( .A1(n89), .A2(n88), .ZN(n93) );
  NAND2_X1 U219 ( .A1(net46455), .A2(net46444), .ZN(net46454) );
  NAND2_X1 U220 ( .A1(n70), .A2(n74), .ZN(n72) );
  NAND2_X1 U221 ( .A1(n44), .A2(n242), .ZN(n239) );
  INV_X1 U222 ( .A(A[0]), .ZN(n242) );
  NAND2_X1 U223 ( .A1(net46444), .A2(net46456), .ZN(n173) );
  NAND2_X1 U224 ( .A1(B[17]), .A2(A[17]), .ZN(n181) );
  NAND2_X1 U225 ( .A1(B[25]), .A2(A[25]), .ZN(n131) );
  OAI211_X1 U226 ( .C1(n214), .C2(n215), .A(n216), .B(n217), .ZN(net46562) );
  AND2_X1 U227 ( .A1(n219), .A2(n220), .ZN(n216) );
  NAND2_X1 U228 ( .A1(n218), .A2(n54), .ZN(n214) );
  OR2_X1 U229 ( .A1(B[17]), .A2(A[17]), .ZN(net46479) );
  OR2_X1 U230 ( .A1(B[26]), .A2(A[26]), .ZN(n126) );
  OR2_X1 U231 ( .A1(B[28]), .A2(A[28]), .ZN(n102) );
  OR2_X1 U232 ( .A1(B[23]), .A2(A[23]), .ZN(n170) );
  OR2_X1 U233 ( .A1(B[16]), .A2(A[16]), .ZN(net46478) );
  OR2_X1 U234 ( .A1(B[21]), .A2(A[21]), .ZN(net46439) );
  INV_X1 U235 ( .A(A[24]), .ZN(n133) );
  OAI21_X1 U236 ( .B1(n123), .B2(n124), .A(n125), .ZN(n122) );
  NAND2_X1 U237 ( .A1(n127), .A2(n126), .ZN(n124) );
  NAND2_X1 U238 ( .A1(n130), .A2(n131), .ZN(n129) );
  OR2_X1 U239 ( .A1(B[11]), .A2(A[11]), .ZN(net46561) );
  OR2_X1 U240 ( .A1(B[6]), .A2(A[6]), .ZN(n60) );
  OR2_X1 U241 ( .A1(B[20]), .A2(A[20]), .ZN(net46443) );
  OR2_X1 U242 ( .A1(B[29]), .A2(A[29]), .ZN(n98) );
  NAND2_X1 U243 ( .A1(n178), .A2(n179), .ZN(net46354) );
  NAND2_X1 U244 ( .A1(n70), .A2(n39), .ZN(n199) );
  OR2_X1 U245 ( .A1(B[30]), .A2(A[30]), .ZN(n89) );
  OR2_X1 U246 ( .A1(B[9]), .A2(A[9]), .ZN(n54) );
  XNOR2_X1 U247 ( .A(n143), .B(n144), .ZN(SUM[27]) );
  NOR2_X1 U248 ( .A1(n224), .A2(n223), .ZN(net46600) );
  OR2_X1 U249 ( .A1(B[7]), .A2(A[7]), .ZN(net46630) );
  OR2_X1 U250 ( .A1(B[19]), .A2(A[19]), .ZN(net46481) );
  OR2_X1 U251 ( .A1(B[4]), .A2(A[4]), .ZN(n74) );
  XNOR2_X1 U252 ( .A(n183), .B(n107), .ZN(SUM[1]) );
  XNOR2_X1 U253 ( .A(n68), .B(n66), .ZN(SUM[5]) );
  XNOR2_X1 U254 ( .A(n103), .B(n79), .ZN(SUM[2]) );
  XNOR2_X1 U255 ( .A(n52), .B(n53), .ZN(SUM[9]) );
  XNOR2_X1 U256 ( .A(n203), .B(net46568), .ZN(SUM[15]) );
  NAND2_X1 U257 ( .A1(net46443), .A2(net46442), .ZN(n177) );
  XNOR2_X1 U258 ( .A(B[31]), .B(A[31]), .ZN(n80) );
  NOR2_X1 U259 ( .A1(n136), .A2(n135), .ZN(n121) );
  NOR2_X1 U260 ( .A1(n135), .A2(n139), .ZN(n138) );
  NAND2_X1 U261 ( .A1(n3), .A2(n57), .ZN(n213) );
  NAND2_X1 U262 ( .A1(B[29]), .A2(A[29]), .ZN(n100) );
  NAND2_X1 U263 ( .A1(B[23]), .A2(A[23]), .ZN(n136) );
  NAND2_X1 U264 ( .A1(B[26]), .A2(A[26]), .ZN(n130) );
  OAI21_X1 U265 ( .B1(n40), .B2(n200), .A(n6), .ZN(n57) );
  OAI21_X1 U266 ( .B1(n69), .B2(n40), .A(n70), .ZN(n66) );
  NAND2_X1 U267 ( .A1(B[5]), .A2(n48), .ZN(n65) );
  XNOR2_X1 U268 ( .A(n177), .B(n176), .ZN(SUM[20]) );
  NAND2_X1 U269 ( .A1(A[11]), .A2(B[11]), .ZN(n219) );
  NOR2_X1 U270 ( .A1(A[11]), .A2(B[11]), .ZN(n224) );
  NAND2_X1 U271 ( .A1(B[27]), .A2(A[27]), .ZN(n125) );
  NAND2_X1 U272 ( .A1(B[4]), .A2(A[4]), .ZN(n70) );
  NAND4_X1 U273 ( .A1(net46303), .A2(A[1]), .A3(n108), .A4(B[1]), .ZN(net46546) );
  NAND2_X1 U274 ( .A1(B[19]), .A2(A[19]), .ZN(net46355) );
  NAND2_X1 U275 ( .A1(B[7]), .A2(n2), .ZN(net46536) );
  OAI22_X1 U276 ( .A1(A[6]), .A2(B[6]), .B1(B[7]), .B2(A[7]), .ZN(n235) );
  NAND2_X1 U277 ( .A1(B[28]), .A2(A[28]), .ZN(n99) );
  OAI211_X1 U278 ( .C1(A[22]), .C2(n13), .A(n170), .B(net46439), .ZN(n140) );
  NAND2_X1 U279 ( .A1(B[18]), .A2(A[18]), .ZN(n182) );
  NAND2_X1 U280 ( .A1(n10), .A2(n4), .ZN(n55) );
  NOR2_X1 U281 ( .A1(B[9]), .A2(A[9]), .ZN(n222) );
  NAND2_X1 U282 ( .A1(B[24]), .A2(A[24]), .ZN(n155) );
  AOI21_X1 U283 ( .B1(n128), .B2(B[24]), .A(n129), .ZN(n123) );
  NAND2_X1 U284 ( .A1(B[10]), .A2(A[10]), .ZN(n220) );
  NOR2_X1 U285 ( .A1(B[10]), .A2(A[10]), .ZN(n223) );
  NAND2_X1 U286 ( .A1(B[30]), .A2(A[30]), .ZN(n88) );
  XNOR2_X1 U287 ( .A(n109), .B(n110), .ZN(SUM[29]) );
  AOI21_X1 U288 ( .B1(n201), .B2(n211), .A(net46588), .ZN(n210) );
  NAND2_X1 U289 ( .A1(B[8]), .A2(A[8]), .ZN(n215) );
  NAND2_X1 U290 ( .A1(net46652), .A2(net46653), .ZN(n202) );
  AOI21_X1 U291 ( .B1(n187), .B2(net46480), .A(n188), .ZN(n185) );
  NAND2_X1 U292 ( .A1(n232), .A2(n215), .ZN(n52) );
  XNOR2_X1 U293 ( .A(n225), .B(n226), .ZN(SUM[11]) );
  NAND2_X1 U294 ( .A1(n227), .A2(n220), .ZN(n225) );
  NAND2_X1 U295 ( .A1(B[16]), .A2(A[16]), .ZN(n194) );
  NAND2_X1 U296 ( .A1(n11), .A2(net52718), .ZN(n201) );
  XNOR2_X1 U297 ( .A(n185), .B(n186), .ZN(SUM[19]) );
  NAND2_X1 U298 ( .A1(B[2]), .A2(A[2]), .ZN(net46301) );
  XNOR2_X1 U299 ( .A(n16), .B(n229), .ZN(SUM[10]) );
  NAND2_X1 U300 ( .A1(n228), .A2(n218), .ZN(n227) );
  NAND2_X1 U301 ( .A1(n47), .A2(n46), .ZN(net46304) );
  NOR2_X1 U302 ( .A1(n47), .A2(n46), .ZN(n241) );
  INV_X1 U303 ( .A(n66), .ZN(n63) );
  XNOR2_X1 U304 ( .A(n72), .B(n73), .ZN(SUM[4]) );
  XNOR2_X1 U305 ( .A(n75), .B(n76), .ZN(SUM[3]) );
  OAI21_X1 U306 ( .B1(n77), .B2(n78), .A(net46301), .ZN(n76) );
  INV_X1 U307 ( .A(n79), .ZN(n77) );
  XNOR2_X1 U308 ( .A(n81), .B(n80), .ZN(SUM[31]) );
  INV_X1 U309 ( .A(n89), .ZN(n86) );
  INV_X1 U310 ( .A(n90), .ZN(n83) );
  XNOR2_X1 U311 ( .A(n94), .B(n93), .ZN(SUM[30]) );
  OAI21_X1 U312 ( .B1(n49), .B2(n9), .A(n95), .ZN(n94) );
  INV_X1 U313 ( .A(n87), .ZN(n96) );
  INV_X1 U314 ( .A(n101), .ZN(n92) );
  INV_X1 U315 ( .A(n99), .ZN(n113) );
  NAND2_X1 U316 ( .A1(n114), .A2(n102), .ZN(n111) );
  INV_X1 U317 ( .A(n91), .ZN(n114) );
  NAND3_X1 U318 ( .A1(n115), .A2(n20), .A3(net46358), .ZN(net46352) );
  XNOR2_X1 U319 ( .A(n117), .B(n116), .ZN(SUM[28]) );
  OAI21_X1 U320 ( .B1(n49), .B2(n91), .A(n118), .ZN(n117) );
  INV_X1 U321 ( .A(n84), .ZN(n118) );
  NOR2_X1 U322 ( .A1(n132), .A2(n133), .ZN(n128) );
  INV_X1 U323 ( .A(n134), .ZN(n132) );
  NAND3_X1 U324 ( .A1(n147), .A2(n145), .A3(n146), .ZN(n143) );
  NAND3_X1 U325 ( .A1(net46321), .A2(net46404), .A3(n148), .ZN(n147) );
  INV_X1 U326 ( .A(net46412), .ZN(net46404) );
  XNOR2_X1 U327 ( .A(n156), .B(n157), .ZN(SUM[26]) );
  OAI21_X1 U328 ( .B1(n49), .B2(n158), .A(n159), .ZN(n157) );
  INV_X1 U329 ( .A(n131), .ZN(n161) );
  NAND2_X1 U330 ( .A1(n45), .A2(n148), .ZN(n158) );
  INV_X1 U331 ( .A(n162), .ZN(n148) );
  XNOR2_X1 U332 ( .A(n163), .B(n164), .ZN(SUM[25]) );
  OAI21_X1 U333 ( .B1(n162), .B2(n49), .A(n165), .ZN(n164) );
  INV_X1 U334 ( .A(n160), .ZN(n165) );
  INV_X1 U335 ( .A(n142), .ZN(n166) );
  INV_X1 U336 ( .A(n167), .ZN(n141) );
  XNOR2_X1 U337 ( .A(n168), .B(n169), .ZN(SUM[24]) );
  OAI21_X1 U338 ( .B1(n49), .B2(n167), .A(n152), .ZN(n169) );
  XNOR2_X1 U339 ( .A(n172), .B(n171), .ZN(SUM[23]) );
  OAI21_X1 U340 ( .B1(n49), .B2(n173), .A(n174), .ZN(n172) );
  INV_X1 U341 ( .A(net46444), .ZN(net46452) );
  INV_X1 U342 ( .A(net46442), .ZN(net46455) );
  XNOR2_X1 U343 ( .A(net46467), .B(n175), .ZN(SUM[21]) );
  OAI21_X1 U344 ( .B1(n49), .B2(net46469), .A(net46442), .ZN(n175) );
  INV_X1 U345 ( .A(net46443), .ZN(net46469) );
  NAND3_X1 U346 ( .A1(n180), .A2(n181), .A3(n182), .ZN(n179) );
  NAND3_X1 U347 ( .A1(A[16]), .A2(net46479), .A3(B[16]), .ZN(n180) );
  INV_X1 U348 ( .A(net46481), .ZN(net46496) );
  INV_X1 U349 ( .A(n182), .ZN(n188) );
  XNOR2_X1 U350 ( .A(n37), .B(n189), .ZN(SUM[18]) );
  INV_X1 U351 ( .A(n181), .ZN(n193) );
  INV_X1 U352 ( .A(n194), .ZN(n192) );
  XNOR2_X1 U353 ( .A(n195), .B(n196), .ZN(SUM[17]) );
  INV_X1 U354 ( .A(net46478), .ZN(net46522) );
  XNOR2_X1 U355 ( .A(n197), .B(net46523), .ZN(SUM[16]) );
  NAND3_X1 U356 ( .A1(n199), .A2(n71), .A3(n198), .ZN(net46488) );
  INV_X1 U357 ( .A(net46556), .ZN(net46571) );
  XNOR2_X1 U358 ( .A(n206), .B(n207), .ZN(SUM[13]) );
  NAND2_X1 U359 ( .A1(n205), .A2(net46579), .ZN(n207) );
  NOR2_X1 U360 ( .A1(n40), .A2(n200), .ZN(n208) );
  NAND3_X1 U361 ( .A1(n218), .A2(n10), .A3(n4), .ZN(n217) );
  NOR2_X1 U362 ( .A1(n221), .A2(n222), .ZN(net46601) );
  INV_X1 U363 ( .A(n58), .ZN(n221) );
  INV_X1 U364 ( .A(n54), .ZN(n231) );
  INV_X1 U365 ( .A(n52), .ZN(n230) );
  NAND2_X1 U366 ( .A1(n233), .A2(n58), .ZN(n232) );
  OAI21_X1 U367 ( .B1(n40), .B2(n200), .A(n6), .ZN(n233) );
  NAND3_X1 U368 ( .A1(n198), .A2(n71), .A3(n234), .ZN(net46626) );
  INV_X1 U369 ( .A(n235), .ZN(n198) );
  NOR2_X1 U370 ( .A1(n19), .A2(n236), .ZN(net46632) );
  INV_X1 U371 ( .A(n60), .ZN(n236) );
  INV_X1 U372 ( .A(n74), .ZN(n69) );
  INV_X1 U373 ( .A(n71), .ZN(n64) );
  NOR2_X1 U374 ( .A1(n240), .A2(n238), .ZN(net46653) );
  NAND2_X1 U375 ( .A1(n43), .A2(A[0]), .ZN(n240) );
  INV_X1 U376 ( .A(n106), .ZN(n238) );
  NOR2_X1 U377 ( .A1(n36), .A2(n241), .ZN(net46652) );
  INV_X1 U378 ( .A(n108), .ZN(n78) );
endmodule


module ALU_N32_DW01_cmp6_5 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428;

  OR2_X1 U1 ( .A1(n375), .A2(B[26]), .ZN(n61) );
  NAND2_X1 U2 ( .A1(A[23]), .A2(n411), .ZN(n64) );
  NAND2_X1 U3 ( .A1(n1), .A2(n2), .ZN(n76) );
  AND2_X1 U4 ( .A1(n10), .A2(n4), .ZN(n1) );
  AND2_X1 U5 ( .A1(n121), .A2(n122), .ZN(n2) );
  AND2_X2 U6 ( .A1(n384), .A2(n72), .ZN(n3) );
  INV_X1 U7 ( .A(n116), .ZN(n4) );
  NAND2_X2 U8 ( .A1(A[20]), .A2(n427), .ZN(n87) );
  AND2_X2 U9 ( .A1(n29), .A2(n364), .ZN(n24) );
  INV_X1 U10 ( .A(A[25]), .ZN(n262) );
  AND2_X1 U11 ( .A1(B[19]), .A2(n20), .ZN(n5) );
  AND2_X1 U12 ( .A1(B[17]), .A2(n242), .ZN(n6) );
  AND3_X1 U13 ( .A1(n24), .A2(n396), .A3(n397), .ZN(n7) );
  AND2_X1 U14 ( .A1(n17), .A2(n232), .ZN(n8) );
  AND2_X1 U15 ( .A1(n267), .A2(n232), .ZN(n9) );
  AND2_X1 U16 ( .A1(n115), .A2(n114), .ZN(n10) );
  AND2_X1 U17 ( .A1(n249), .A2(n247), .ZN(n11) );
  AND2_X1 U18 ( .A1(n236), .A2(n235), .ZN(n12) );
  BUF_X1 U19 ( .A(n92), .Z(n13) );
  NOR3_X1 U20 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n220) );
  NOR2_X1 U21 ( .A1(n265), .A2(n266), .ZN(n14) );
  AND4_X1 U22 ( .A1(n17), .A2(n263), .A3(n232), .A4(n24), .ZN(n15) );
  NOR2_X1 U23 ( .A1(n33), .A2(n261), .ZN(n16) );
  AND2_X2 U24 ( .A1(n86), .A2(n61), .ZN(n17) );
  NAND2_X1 U25 ( .A1(B[10]), .A2(n329), .ZN(n284) );
  NAND2_X2 U26 ( .A1(A[24]), .A2(n405), .ZN(n63) );
  INV_X1 U27 ( .A(n85), .ZN(n18) );
  AND2_X2 U28 ( .A1(B[31]), .A2(n131), .ZN(n19) );
  INV_X2 U29 ( .A(n19), .ZN(n232) );
  INV_X1 U30 ( .A(n24), .ZN(n33) );
  NAND2_X2 U31 ( .A1(n407), .A2(A[18]), .ZN(n93) );
  OR2_X2 U32 ( .A1(B[19]), .A2(n20), .ZN(n120) );
  INV_X1 U33 ( .A(A[19]), .ZN(n20) );
  AND2_X1 U34 ( .A1(A[19]), .A2(n404), .ZN(n21) );
  BUF_X1 U35 ( .A(n123), .Z(n22) );
  CLKBUF_X1 U36 ( .A(B[18]), .Z(n23) );
  NAND3_X1 U37 ( .A1(n248), .A2(n231), .A3(n8), .ZN(n291) );
  NAND2_X1 U38 ( .A1(n75), .A2(n362), .ZN(n25) );
  NAND2_X1 U39 ( .A1(n362), .A2(n75), .ZN(n26) );
  NAND2_X1 U40 ( .A1(n75), .A2(n362), .ZN(n132) );
  AND2_X1 U41 ( .A1(n258), .A2(n93), .ZN(n27) );
  NAND3_X1 U42 ( .A1(n238), .A2(n237), .A3(n12), .ZN(n224) );
  NAND2_X1 U43 ( .A1(n86), .A2(n61), .ZN(n28) );
  NOR2_X1 U44 ( .A1(n18), .A2(n417), .ZN(n29) );
  NOR2_X1 U45 ( .A1(n18), .A2(n417), .ZN(n414) );
  NAND3_X1 U46 ( .A1(n248), .A2(n369), .A3(n11), .ZN(n246) );
  NAND2_X1 U47 ( .A1(n252), .A2(n58), .ZN(n30) );
  INV_X1 U48 ( .A(n87), .ZN(n31) );
  NAND3_X1 U49 ( .A1(n24), .A2(n268), .A3(n9), .ZN(n266) );
  NAND2_X1 U50 ( .A1(n414), .A2(n364), .ZN(n32) );
  INV_X1 U51 ( .A(n88), .ZN(n34) );
  AND2_X2 U52 ( .A1(n398), .A2(n87), .ZN(n35) );
  NOR2_X1 U53 ( .A1(n132), .A2(n19), .ZN(n249) );
  OAI21_X1 U54 ( .B1(n188), .B2(n189), .A(n190), .ZN(n176) );
  AOI21_X1 U55 ( .B1(n191), .B2(n192), .A(n111), .ZN(n190) );
  AOI21_X1 U56 ( .B1(n378), .B2(n379), .A(n380), .ZN(n354) );
  NAND2_X1 U57 ( .A1(n381), .A2(n382), .ZN(n380) );
  NOR2_X1 U58 ( .A1(n390), .A2(n389), .ZN(n378) );
  NOR2_X1 U59 ( .A1(n386), .A2(n387), .ZN(n379) );
  AOI21_X1 U60 ( .B1(n394), .B2(n395), .A(n7), .ZN(n353) );
  NOR2_X1 U61 ( .A1(n412), .A2(n413), .ZN(n394) );
  NOR2_X1 U62 ( .A1(n386), .A2(n400), .ZN(n395) );
  NOR2_X1 U63 ( .A1(n158), .A2(n170), .ZN(n192) );
  NAND2_X1 U64 ( .A1(n224), .A2(n225), .ZN(n223) );
  OAI211_X1 U65 ( .C1(n243), .C2(n244), .A(n245), .B(n246), .ZN(n222) );
  NOR2_X1 U66 ( .A1(n76), .A2(n77), .ZN(n41) );
  NOR2_X1 U67 ( .A1(n47), .A2(n48), .ZN(n46) );
  NOR2_X1 U68 ( .A1(n250), .A2(n251), .ZN(n369) );
  NOR2_X1 U69 ( .A1(n145), .A2(n146), .ZN(n144) );
  NAND4_X1 U70 ( .A1(n297), .A2(n296), .A3(n295), .A4(n298), .ZN(n218) );
  NOR2_X1 U71 ( .A1(n34), .A2(n351), .ZN(n295) );
  NOR2_X1 U72 ( .A1(n299), .A2(n300), .ZN(n298) );
  INV_X1 U73 ( .A(n305), .ZN(n304) );
  OR2_X1 U74 ( .A1(n30), .A2(n26), .ZN(n399) );
  NOR2_X1 U75 ( .A1(n276), .A2(n277), .ZN(n275) );
  NOR2_X1 U76 ( .A1(n147), .A2(n148), .ZN(n142) );
  INV_X1 U77 ( .A(n113), .ZN(n292) );
  NAND2_X1 U78 ( .A1(n69), .A2(n62), .ZN(n417) );
  NAND2_X1 U79 ( .A1(n284), .A2(n215), .ZN(n145) );
  NAND2_X1 U80 ( .A1(n205), .A2(n281), .ZN(n170) );
  INV_X1 U81 ( .A(n99), .ZN(n370) );
  INV_X1 U82 ( .A(n74), .ZN(n363) );
  NAND4_X1 U83 ( .A1(n3), .A2(n69), .A3(n361), .A4(n232), .ZN(n360) );
  INV_X1 U84 ( .A(n362), .ZN(n361) );
  NAND4_X1 U85 ( .A1(n17), .A2(n388), .A3(n36), .A4(n232), .ZN(n261) );
  NAND2_X1 U86 ( .A1(n106), .A2(n174), .ZN(n305) );
  NAND2_X1 U87 ( .A1(n232), .A2(n385), .ZN(n381) );
  INV_X1 U88 ( .A(n70), .ZN(n385) );
  NAND2_X1 U89 ( .A1(n383), .A2(n232), .ZN(n382) );
  INV_X1 U90 ( .A(n384), .ZN(n383) );
  NAND2_X1 U91 ( .A1(n187), .A2(n287), .ZN(n148) );
  NAND2_X1 U92 ( .A1(n318), .A2(n196), .ZN(n146) );
  AND2_X1 U93 ( .A1(n64), .A2(n120), .ZN(n259) );
  NOR2_X1 U94 ( .A1(n250), .A2(n25), .ZN(n260) );
  INV_X1 U95 ( .A(n293), .ZN(n391) );
  NAND2_X1 U96 ( .A1(n99), .A2(n57), .ZN(n98) );
  NOR2_X1 U97 ( .A1(n100), .A2(n101), .ZN(n97) );
  NOR2_X1 U98 ( .A1(n103), .A2(n104), .ZN(n96) );
  NOR3_X1 U99 ( .A1(n356), .A2(n357), .A3(n358), .ZN(n355) );
  NAND2_X1 U100 ( .A1(n359), .A2(n360), .ZN(n358) );
  NOR2_X1 U101 ( .A1(n366), .A2(n367), .ZN(n357) );
  AOI21_X1 U102 ( .B1(n313), .B2(n314), .A(n315), .ZN(n297) );
  AND3_X1 U103 ( .A1(n320), .A2(n183), .A3(n287), .ZN(n314) );
  NOR2_X1 U104 ( .A1(n322), .A2(n305), .ZN(n313) );
  NOR2_X1 U105 ( .A1(n316), .A2(n317), .ZN(n315) );
  OAI211_X1 U106 ( .C1(n278), .C2(n279), .A(n119), .B(n280), .ZN(n276) );
  NAND2_X1 U107 ( .A1(n288), .A2(n183), .ZN(n278) );
  NAND4_X1 U108 ( .A1(n281), .A2(n282), .A3(n283), .A4(n284), .ZN(n280) );
  NAND4_X1 U109 ( .A1(n287), .A2(n284), .A3(n281), .A4(n282), .ZN(n279) );
  AND3_X1 U110 ( .A1(n6), .A2(n63), .A3(n64), .ZN(n235) );
  NOR2_X1 U111 ( .A1(n123), .A2(n241), .ZN(n236) );
  NOR2_X1 U112 ( .A1(n19), .A2(n240), .ZN(n237) );
  INV_X1 U113 ( .A(n212), .ZN(n310) );
  NAND4_X1 U114 ( .A1(n281), .A2(n287), .A3(n183), .A4(n282), .ZN(n317) );
  NAND4_X1 U115 ( .A1(n281), .A2(n284), .A3(n175), .A4(n318), .ZN(n322) );
  NAND4_X1 U116 ( .A1(n67), .A2(n129), .A3(n74), .A4(n130), .ZN(n47) );
  NAND4_X1 U117 ( .A1(n64), .A2(n91), .A3(n88), .A4(n27), .ZN(n386) );
  NAND4_X1 U118 ( .A1(n284), .A2(n175), .A3(n318), .A4(n146), .ZN(n316) );
  OAI211_X1 U119 ( .C1(n301), .C2(n302), .A(n64), .B(n303), .ZN(n300) );
  NAND4_X1 U120 ( .A1(n145), .A2(n284), .A3(n281), .A4(n304), .ZN(n303) );
  OAI21_X1 U121 ( .B1(n167), .B2(n168), .A(n91), .ZN(n137) );
  INV_X1 U122 ( .A(n128), .ZN(n401) );
  INV_X1 U123 ( .A(n26), .ZN(n388) );
  NAND2_X1 U124 ( .A1(n258), .A2(n93), .ZN(n123) );
  NOR2_X1 U125 ( .A1(n54), .A2(n64), .ZN(n59) );
  OAI21_X1 U126 ( .B1(n139), .B2(n140), .A(n141), .ZN(n138) );
  OAI211_X1 U127 ( .C1(n149), .C2(n150), .A(n151), .B(n152), .ZN(n139) );
  OAI21_X1 U128 ( .B1(n160), .B2(n161), .A(n162), .ZN(n150) );
  NOR2_X1 U129 ( .A1(n145), .A2(n193), .ZN(n191) );
  NOR2_X1 U130 ( .A1(n153), .A2(n154), .ZN(n152) );
  NAND2_X1 U131 ( .A1(n155), .A2(n156), .ZN(n154) );
  NAND4_X1 U132 ( .A1(n253), .A2(n24), .A3(n50), .A4(n254), .ZN(n245) );
  NOR2_X1 U133 ( .A1(n28), .A2(n57), .ZN(n253) );
  NOR2_X1 U134 ( .A1(n250), .A2(n19), .ZN(n254) );
  NAND2_X1 U135 ( .A1(n88), .A2(n120), .ZN(n241) );
  NOR2_X1 U136 ( .A1(n28), .A2(n252), .ZN(n247) );
  NOR2_X1 U137 ( .A1(n54), .A2(n55), .ZN(n53) );
  NAND2_X1 U138 ( .A1(n91), .A2(n120), .ZN(n272) );
  NOR3_X1 U139 ( .A1(n19), .A2(n398), .A3(n28), .ZN(n397) );
  NOR2_X1 U140 ( .A1(n233), .A2(n399), .ZN(n396) );
  NAND4_X1 U141 ( .A1(n17), .A2(n114), .A3(n232), .A4(n24), .ZN(n413) );
  AND4_X1 U142 ( .A1(n200), .A2(n88), .A3(n201), .A4(n202), .ZN(n134) );
  NOR2_X1 U143 ( .A1(n137), .A2(n138), .ZN(n136) );
  NOR2_X1 U144 ( .A1(n176), .A2(n177), .ZN(n135) );
  NAND2_X1 U145 ( .A1(n93), .A2(n102), .ZN(n100) );
  NAND2_X1 U146 ( .A1(n269), .A2(n92), .ZN(n94) );
  NOR2_X1 U147 ( .A1(n170), .A2(n186), .ZN(n185) );
  NAND2_X1 U148 ( .A1(n174), .A2(n183), .ZN(n186) );
  NOR2_X1 U149 ( .A1(n25), .A2(n273), .ZN(n270) );
  NOR2_X1 U150 ( .A1(n34), .A2(n272), .ZN(n271) );
  NAND2_X1 U151 ( .A1(n64), .A2(n63), .ZN(n273) );
  NAND2_X1 U152 ( .A1(n13), .A2(n204), .ZN(n351) );
  NOR2_X1 U153 ( .A1(n182), .A2(n145), .ZN(n181) );
  NOR2_X1 U154 ( .A1(n19), .A2(n230), .ZN(n227) );
  OAI21_X1 U155 ( .B1(n117), .B2(n118), .A(n119), .ZN(n116) );
  NOR2_X1 U156 ( .A1(n345), .A2(n305), .ZN(n323) );
  NAND2_X1 U157 ( .A1(n84), .A2(n85), .ZN(n49) );
  NOR2_X1 U158 ( .A1(n233), .A2(n234), .ZN(n226) );
  NAND2_X1 U159 ( .A1(n50), .A2(n5), .ZN(n234) );
  NOR2_X1 U160 ( .A1(n31), .A2(n203), .ZN(n202) );
  NAND4_X1 U161 ( .A1(n204), .A2(n205), .A3(n102), .A4(n93), .ZN(n203) );
  NOR2_X1 U162 ( .A1(n110), .A2(n103), .ZN(n109) );
  NOR2_X1 U163 ( .A1(n81), .A2(n82), .ZN(n80) );
  NOR2_X1 U164 ( .A1(n89), .A2(n90), .ZN(n81) );
  NOR2_X1 U165 ( .A1(n145), .A2(n187), .ZN(n184) );
  AND2_X1 U166 ( .A1(n232), .A2(n17), .ZN(n257) );
  OAI21_X1 U167 ( .B1(n65), .B2(n66), .A(n67), .ZN(n43) );
  AND3_X1 U168 ( .A1(n113), .A2(n102), .A3(n93), .ZN(n107) );
  OR2_X1 U169 ( .A1(n372), .A2(n129), .ZN(n373) );
  NAND2_X1 U170 ( .A1(n51), .A2(n52), .ZN(n45) );
  NOR2_X1 U171 ( .A1(n59), .A2(n60), .ZN(n51) );
  NOR2_X1 U172 ( .A1(n18), .A2(n53), .ZN(n52) );
  OAI21_X1 U173 ( .B1(n164), .B2(n165), .A(n166), .ZN(n149) );
  OAI21_X1 U174 ( .B1(A[1]), .B2(n38), .A(A[0]), .ZN(n165) );
  NAND2_X1 U175 ( .A1(n163), .A2(n37), .ZN(n164) );
  NAND2_X1 U176 ( .A1(n293), .A2(n102), .ZN(n113) );
  NOR2_X1 U177 ( .A1(n209), .A2(n146), .ZN(n206) );
  NOR2_X1 U178 ( .A1(n153), .A2(n199), .ZN(n208) );
  NOR2_X1 U179 ( .A1(n170), .A2(n145), .ZN(n207) );
  NOR2_X1 U180 ( .A1(n343), .A2(n344), .ZN(n340) );
  NOR2_X1 U181 ( .A1(A[0]), .A2(n37), .ZN(n343) );
  NAND2_X1 U182 ( .A1(A[1]), .A2(n38), .ZN(n161) );
  OAI21_X1 U183 ( .B1(n333), .B2(n334), .A(n335), .ZN(n324) );
  NAND2_X1 U184 ( .A1(n156), .A2(n163), .ZN(n334) );
  AND2_X1 U185 ( .A1(n171), .A2(n162), .ZN(n335) );
  NOR2_X1 U186 ( .A1(n340), .A2(n341), .ZN(n333) );
  NOR2_X1 U187 ( .A1(n153), .A2(n173), .ZN(n172) );
  NAND2_X1 U188 ( .A1(n174), .A2(n159), .ZN(n173) );
  NOR2_X1 U189 ( .A1(n153), .A2(n199), .ZN(n197) );
  NAND2_X1 U190 ( .A1(n174), .A2(n175), .ZN(n199) );
  NOR2_X1 U191 ( .A1(n146), .A2(n171), .ZN(n169) );
  NOR2_X1 U192 ( .A1(n148), .A2(n186), .ZN(n180) );
  NOR2_X1 U193 ( .A1(n326), .A2(n327), .ZN(n325) );
  NAND2_X1 U194 ( .A1(n284), .A2(n175), .ZN(n327) );
  NOR2_X1 U195 ( .A1(n210), .A2(n211), .ZN(n200) );
  NOR2_X1 U196 ( .A1(n170), .A2(n213), .ZN(n210) );
  NOR2_X1 U197 ( .A1(n170), .A2(n212), .ZN(n211) );
  NAND2_X1 U198 ( .A1(n342), .A2(n166), .ZN(n341) );
  NAND2_X1 U199 ( .A1(A[1]), .A2(n38), .ZN(n342) );
  INV_X1 U200 ( .A(n182), .ZN(n288) );
  INV_X1 U201 ( .A(n193), .ZN(n283) );
  INV_X1 U202 ( .A(n209), .ZN(n320) );
  INV_X1 U203 ( .A(A[31]), .ZN(n131) );
  INV_X1 U204 ( .A(B[17]), .ZN(n410) );
  NAND2_X1 U205 ( .A1(B[11]), .A2(n346), .ZN(n174) );
  NAND2_X1 U206 ( .A1(A[16]), .A2(n425), .ZN(n92) );
  NOR2_X1 U207 ( .A1(n25), .A2(n286), .ZN(n263) );
  NAND2_X1 U208 ( .A1(B[8]), .A2(n350), .ZN(n287) );
  NAND2_X1 U209 ( .A1(A[29]), .A2(n419), .ZN(n69) );
  INV_X1 U210 ( .A(B[12]), .ZN(n312) );
  INV_X1 U211 ( .A(A[28]), .ZN(n424) );
  INV_X1 U212 ( .A(A[17]), .ZN(n242) );
  NAND2_X1 U213 ( .A1(n423), .A2(A[28]), .ZN(n75) );
  INV_X1 U214 ( .A(A[23]), .ZN(n255) );
  INV_X1 U215 ( .A(B[6]), .ZN(n319) );
  NAND2_X1 U216 ( .A1(A[27]), .A2(n420), .ZN(n85) );
  NAND2_X1 U217 ( .A1(B[13]), .A2(n347), .ZN(n106) );
  INV_X1 U218 ( .A(A[18]), .ZN(n408) );
  NAND2_X1 U219 ( .A1(n286), .A2(n63), .ZN(n54) );
  NAND2_X1 U220 ( .A1(n120), .A2(n402), .ZN(n103) );
  INV_X1 U221 ( .A(B[10]), .ZN(n306) );
  NAND2_X1 U222 ( .A1(B[6]), .A2(n332), .ZN(n318) );
  INV_X1 U223 ( .A(A[20]), .ZN(n428) );
  INV_X1 U224 ( .A(A[22]), .ZN(n422) );
  INV_X1 U225 ( .A(A[24]), .ZN(n264) );
  INV_X1 U226 ( .A(A[16]), .ZN(n426) );
  INV_X1 U227 ( .A(A[30]), .ZN(n416) );
  INV_X1 U228 ( .A(A[26]), .ZN(n375) );
  INV_X1 U229 ( .A(B[14]), .ZN(n294) );
  INV_X1 U230 ( .A(B[11]), .ZN(n311) );
  INV_X1 U231 ( .A(A[29]), .ZN(n365) );
  INV_X1 U232 ( .A(B[5]), .ZN(n321) );
  INV_X1 U233 ( .A(A[27]), .ZN(n374) );
  NAND2_X1 U234 ( .A1(A[2]), .A2(n39), .ZN(n166) );
  NAND2_X1 U235 ( .A1(B[5]), .A2(n330), .ZN(n159) );
  INV_X1 U236 ( .A(B[7]), .ZN(n289) );
  INV_X1 U237 ( .A(B[8]), .ZN(n307) );
  INV_X1 U238 ( .A(B[13]), .ZN(n352) );
  INV_X1 U239 ( .A(A[21]), .ZN(n371) );
  NAND2_X1 U240 ( .A1(B[14]), .A2(n393), .ZN(n293) );
  AND2_X1 U241 ( .A1(B[25]), .A2(n262), .ZN(n36) );
  INV_X1 U242 ( .A(A[2]), .ZN(n338) );
  NAND2_X1 U243 ( .A1(B[7]), .A2(n328), .ZN(n175) );
  OR2_X1 U244 ( .A1(B[31]), .A2(n131), .ZN(n67) );
  AOI21_X1 U245 ( .B1(n41), .B2(n40), .A(n42), .ZN(LE) );
  NAND2_X1 U246 ( .A1(A[25]), .A2(n418), .ZN(n62) );
  INV_X1 U247 ( .A(B[25]), .ZN(n418) );
  NAND2_X1 U248 ( .A1(n384), .A2(n72), .ZN(n68) );
  NAND2_X1 U249 ( .A1(n252), .A2(n58), .ZN(n133) );
  NAND2_X1 U250 ( .A1(A[22]), .A2(n421), .ZN(n58) );
  NAND2_X1 U251 ( .A1(n274), .A2(n275), .ZN(n219) );
  NAND2_X1 U252 ( .A1(B[4]), .A2(n331), .ZN(n155) );
  INV_X1 U253 ( .A(B[4]), .ZN(n337) );
  XNOR2_X1 U254 ( .A(B[31]), .B(A[31]), .ZN(n70) );
  NOR2_X1 U255 ( .A1(n229), .A2(n258), .ZN(n256) );
  NOR2_X1 U256 ( .A1(n269), .A2(n229), .ZN(n268) );
  NOR2_X1 U257 ( .A1(n25), .A2(n30), .ZN(n114) );
  NOR2_X1 U258 ( .A1(n133), .A2(n28), .ZN(n267) );
  NOR2_X1 U259 ( .A1(n30), .A2(n25), .ZN(n368) );
  NAND2_X1 U260 ( .A1(B[29]), .A2(n365), .ZN(n74) );
  INV_X1 U261 ( .A(B[29]), .ZN(n419) );
  OAI21_X1 U262 ( .B1(n372), .B2(n86), .A(n373), .ZN(n356) );
  NAND2_X1 U263 ( .A1(A[30]), .A2(n415), .ZN(n72) );
  NAND2_X1 U264 ( .A1(B[23]), .A2(n255), .ZN(n57) );
  INV_X1 U265 ( .A(B[23]), .ZN(n411) );
  NAND4_X1 U266 ( .A1(n107), .A2(n87), .A3(n108), .A4(n109), .ZN(n78) );
  NAND2_X1 U267 ( .A1(n88), .A2(n87), .ZN(n101) );
  NAND2_X1 U268 ( .A1(B[26]), .A2(n375), .ZN(n86) );
  NAND2_X1 U269 ( .A1(A[5]), .A2(n321), .ZN(n209) );
  INV_X1 U270 ( .A(A[5]), .ZN(n330) );
  NAND2_X1 U271 ( .A1(A[3]), .A2(n336), .ZN(n162) );
  INV_X1 U272 ( .A(A[3]), .ZN(n339) );
  NAND2_X1 U273 ( .A1(A[11]), .A2(n311), .ZN(n212) );
  INV_X1 U274 ( .A(A[11]), .ZN(n346) );
  NAND2_X1 U275 ( .A1(A[12]), .A2(n312), .ZN(n205) );
  INV_X1 U276 ( .A(A[12]), .ZN(n348) );
  OAI211_X1 U277 ( .C1(n35), .C2(n101), .A(n83), .B(n49), .ZN(n82) );
  NAND2_X1 U278 ( .A1(n35), .A2(n292), .ZN(n290) );
  NAND4_X1 U279 ( .A1(n392), .A2(n391), .A3(n35), .A4(n24), .ZN(n390) );
  NAND2_X1 U280 ( .A1(n35), .A2(n392), .ZN(n412) );
  OAI21_X1 U281 ( .B1(n68), .B2(n69), .A(n70), .ZN(n66) );
  OAI21_X1 U282 ( .B1(n68), .B2(n71), .A(n72), .ZN(n65) );
  NOR2_X1 U283 ( .A1(n47), .A2(n68), .ZN(n115) );
  INV_X1 U284 ( .A(n68), .ZN(n364) );
  INV_X1 U285 ( .A(A[15]), .ZN(n406) );
  NAND2_X1 U286 ( .A1(A[15]), .A2(n403), .ZN(n402) );
  NAND2_X1 U287 ( .A1(B[27]), .A2(n374), .ZN(n129) );
  INV_X1 U288 ( .A(B[27]), .ZN(n420) );
  NAND2_X1 U289 ( .A1(A[4]), .A2(n337), .ZN(n171) );
  INV_X1 U290 ( .A(A[4]), .ZN(n331) );
  NAND2_X1 U291 ( .A1(n231), .A2(n17), .ZN(n230) );
  NAND2_X1 U292 ( .A1(n388), .A2(n231), .ZN(n240) );
  NAND4_X1 U293 ( .A1(n259), .A2(n88), .A3(n231), .A4(n260), .ZN(n243) );
  NAND2_X1 U294 ( .A1(A[9]), .A2(n285), .ZN(n193) );
  INV_X1 U295 ( .A(A[9]), .ZN(n349) );
  NOR2_X1 U296 ( .A1(A[1]), .A2(n38), .ZN(n344) );
  INV_X1 U297 ( .A(B[19]), .ZN(n404) );
  NAND2_X1 U298 ( .A1(A[6]), .A2(n319), .ZN(n196) );
  INV_X1 U299 ( .A(A[6]), .ZN(n332) );
  NAND2_X1 U300 ( .A1(A[14]), .A2(n294), .ZN(n102) );
  INV_X1 U301 ( .A(A[14]), .ZN(n393) );
  NAND2_X1 U302 ( .A1(A[13]), .A2(n352), .ZN(n204) );
  INV_X1 U303 ( .A(A[13]), .ZN(n347) );
  NAND2_X1 U304 ( .A1(A[7]), .A2(n289), .ZN(n182) );
  INV_X1 U305 ( .A(A[7]), .ZN(n328) );
  NAND2_X1 U306 ( .A1(B[20]), .A2(n428), .ZN(n398) );
  INV_X1 U307 ( .A(B[20]), .ZN(n427) );
  NAND2_X1 U308 ( .A1(B[28]), .A2(n424), .ZN(n362) );
  INV_X1 U309 ( .A(B[28]), .ZN(n423) );
  NAND2_X1 U310 ( .A1(B[21]), .A2(n371), .ZN(n99) );
  INV_X1 U311 ( .A(B[21]), .ZN(n409) );
  NAND2_X1 U312 ( .A1(B[15]), .A2(n406), .ZN(n128) );
  INV_X1 U313 ( .A(B[15]), .ZN(n403) );
  NAND2_X1 U314 ( .A1(B[22]), .A2(n422), .ZN(n252) );
  INV_X1 U315 ( .A(B[22]), .ZN(n421) );
  NAND2_X1 U316 ( .A1(n23), .A2(n408), .ZN(n258) );
  INV_X1 U317 ( .A(B[18]), .ZN(n407) );
  INV_X1 U318 ( .A(B[9]), .ZN(n285) );
  NAND2_X1 U319 ( .A1(B[9]), .A2(n349), .ZN(n183) );
  NAND2_X1 U320 ( .A1(B[24]), .A2(n264), .ZN(n286) );
  INV_X1 U321 ( .A(B[24]), .ZN(n405) );
  NAND2_X1 U322 ( .A1(A[10]), .A2(n306), .ZN(n215) );
  INV_X1 U323 ( .A(A[10]), .ZN(n329) );
  NOR2_X1 U324 ( .A1(n291), .A2(n290), .ZN(n274) );
  NAND4_X1 U325 ( .A1(n232), .A2(n50), .A3(n376), .A4(n3), .ZN(n372) );
  NAND2_X1 U326 ( .A1(B[30]), .A2(n416), .ZN(n384) );
  INV_X1 U327 ( .A(B[30]), .ZN(n415) );
  NAND2_X1 U328 ( .A1(A[8]), .A2(n307), .ZN(n187) );
  INV_X1 U329 ( .A(A[8]), .ZN(n350) );
  NAND2_X1 U330 ( .A1(B[16]), .A2(n426), .ZN(n269) );
  INV_X1 U331 ( .A(B[16]), .ZN(n425) );
  NOR2_X1 U332 ( .A1(n222), .A2(n223), .ZN(n221) );
  NAND2_X1 U333 ( .A1(B[2]), .A2(n338), .ZN(n163) );
  NAND2_X1 U334 ( .A1(B[3]), .A2(n339), .ZN(n156) );
  INV_X1 U335 ( .A(B[3]), .ZN(n336) );
  NOR2_X1 U336 ( .A1(n217), .A2(n216), .ZN(GE) );
  OAI211_X1 U337 ( .C1(n219), .C2(n218), .A(n221), .B(n220), .ZN(n217) );
  NOR2_X1 U338 ( .A1(n32), .A2(n229), .ZN(n228) );
  INV_X1 U339 ( .A(n32), .ZN(n248) );
  NOR2_X1 U340 ( .A1(n32), .A2(n239), .ZN(n238) );
  NAND2_X1 U341 ( .A1(n35), .A2(n17), .ZN(n239) );
  NAND2_X1 U342 ( .A1(n398), .A2(n87), .ZN(n229) );
  INV_X1 U343 ( .A(B[0]), .ZN(n37) );
  INV_X1 U344 ( .A(B[1]), .ZN(n38) );
  INV_X1 U345 ( .A(B[2]), .ZN(n39) );
  NAND2_X1 U346 ( .A1(n43), .A2(n44), .ZN(n42) );
  NAND2_X1 U347 ( .A1(n45), .A2(n46), .ZN(n44) );
  NAND3_X1 U348 ( .A1(n49), .A2(n3), .A3(n388), .ZN(n48) );
  NAND2_X1 U349 ( .A1(n56), .A2(n57), .ZN(n55) );
  INV_X1 U350 ( .A(n58), .ZN(n56) );
  NAND3_X1 U351 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n60) );
  NAND2_X1 U352 ( .A1(n73), .A2(n74), .ZN(n71) );
  INV_X1 U353 ( .A(n75), .ZN(n73) );
  NAND3_X1 U354 ( .A1(n80), .A2(n79), .A3(n78), .ZN(n77) );
  INV_X1 U355 ( .A(n86), .ZN(n84) );
  NAND3_X1 U356 ( .A1(n5), .A2(n87), .A3(n88), .ZN(n83) );
  NAND3_X1 U357 ( .A1(n91), .A2(n92), .A3(n88), .ZN(n90) );
  NAND3_X1 U358 ( .A1(n93), .A2(n94), .A3(n95), .ZN(n89) );
  NOR2_X1 U359 ( .A1(n31), .A2(n21), .ZN(n95) );
  AOI21_X1 U360 ( .B1(n96), .B2(n97), .A(n98), .ZN(n79) );
  NAND3_X1 U361 ( .A1(n91), .A2(n105), .A3(n92), .ZN(n104) );
  INV_X1 U362 ( .A(n106), .ZN(n105) );
  NOR2_X1 U363 ( .A1(n111), .A2(n34), .ZN(n108) );
  NAND2_X1 U364 ( .A1(n6), .A2(n88), .ZN(n118) );
  NAND3_X1 U365 ( .A1(n120), .A2(n93), .A3(n87), .ZN(n117) );
  NAND3_X1 U366 ( .A1(n127), .A2(n22), .A3(n124), .ZN(n122) );
  NOR2_X1 U367 ( .A1(n21), .A2(n112), .ZN(n124) );
  NAND4_X1 U368 ( .A1(n126), .A2(n13), .A3(n127), .A4(n124), .ZN(n121) );
  NOR2_X1 U369 ( .A1(n125), .A2(n31), .ZN(n127) );
  INV_X1 U370 ( .A(n93), .ZN(n125) );
  NOR2_X1 U371 ( .A1(n128), .A2(n110), .ZN(n126) );
  INV_X1 U372 ( .A(n91), .ZN(n110) );
  NAND3_X1 U373 ( .A1(n36), .A2(n61), .A3(n85), .ZN(n130) );
  NAND3_X1 U374 ( .A1(n134), .A2(n135), .A3(n136), .ZN(n40) );
  NAND3_X1 U375 ( .A1(n142), .A2(n143), .A3(n144), .ZN(n140) );
  NOR2_X1 U376 ( .A1(n157), .A2(n158), .ZN(n151) );
  INV_X1 U377 ( .A(n159), .ZN(n157) );
  INV_X1 U378 ( .A(n163), .ZN(n160) );
  NAND2_X1 U379 ( .A1(n169), .A2(n207), .ZN(n168) );
  NAND2_X1 U380 ( .A1(n142), .A2(n172), .ZN(n167) );
  INV_X1 U381 ( .A(n175), .ZN(n147) );
  NAND2_X1 U382 ( .A1(n178), .A2(n179), .ZN(n177) );
  NAND3_X1 U383 ( .A1(n180), .A2(n143), .A3(n181), .ZN(n179) );
  NAND2_X1 U384 ( .A1(n184), .A2(n185), .ZN(n178) );
  INV_X1 U385 ( .A(n92), .ZN(n111) );
  INV_X1 U386 ( .A(n174), .ZN(n158) );
  NAND3_X1 U387 ( .A1(n194), .A2(n195), .A3(n143), .ZN(n189) );
  INV_X1 U388 ( .A(n170), .ZN(n143) );
  INV_X1 U389 ( .A(n196), .ZN(n195) );
  INV_X1 U390 ( .A(n145), .ZN(n194) );
  NAND2_X1 U391 ( .A1(n197), .A2(n198), .ZN(n188) );
  NAND4_X1 U392 ( .A1(n206), .A2(n207), .A3(n208), .A4(n198), .ZN(n201) );
  INV_X1 U393 ( .A(n148), .ZN(n198) );
  INV_X1 U394 ( .A(n183), .ZN(n153) );
  NAND2_X1 U395 ( .A1(n214), .A2(n174), .ZN(n213) );
  INV_X1 U396 ( .A(n215), .ZN(n214) );
  NAND3_X1 U397 ( .A1(n227), .A2(n226), .A3(n228), .ZN(n225) );
  NAND3_X1 U398 ( .A1(n63), .A2(n88), .A3(n64), .ZN(n233) );
  NAND3_X1 U399 ( .A1(n24), .A2(n256), .A3(n257), .ZN(n244) );
  NAND3_X1 U400 ( .A1(n27), .A2(n270), .A3(n271), .ZN(n265) );
  NAND3_X1 U401 ( .A1(n388), .A2(n27), .A3(n141), .ZN(n277) );
  INV_X1 U402 ( .A(n54), .ZN(n119) );
  NAND3_X1 U403 ( .A1(n183), .A2(n287), .A3(n304), .ZN(n302) );
  NAND3_X1 U404 ( .A1(n284), .A2(n281), .A3(n148), .ZN(n301) );
  NAND3_X1 U405 ( .A1(n308), .A2(n309), .A3(n91), .ZN(n299) );
  NAND3_X1 U406 ( .A1(n281), .A2(n310), .A3(n106), .ZN(n309) );
  NAND3_X1 U407 ( .A1(n106), .A2(n281), .A3(n170), .ZN(n308) );
  INV_X1 U408 ( .A(n305), .ZN(n282) );
  NAND3_X1 U409 ( .A1(n323), .A2(n324), .A3(n325), .ZN(n296) );
  NAND3_X1 U410 ( .A1(n318), .A2(n155), .A3(n159), .ZN(n326) );
  NAND3_X1 U411 ( .A1(n287), .A2(n183), .A3(n281), .ZN(n345) );
  NAND2_X2 U412 ( .A1(B[12]), .A2(n348), .ZN(n281) );
  INV_X1 U413 ( .A(n88), .ZN(n112) );
  NAND3_X1 U414 ( .A1(n353), .A2(n354), .A3(n355), .ZN(n216) );
  NAND3_X1 U415 ( .A1(n363), .A2(n3), .A3(n232), .ZN(n359) );
  NAND3_X1 U416 ( .A1(n368), .A2(n369), .A3(n24), .ZN(n367) );
  INV_X1 U417 ( .A(n64), .ZN(n251) );
  INV_X1 U418 ( .A(n63), .ZN(n250) );
  NAND3_X1 U419 ( .A1(n17), .A2(n370), .A3(n232), .ZN(n366) );
  NOR2_X1 U420 ( .A1(n18), .A2(n377), .ZN(n376) );
  INV_X1 U421 ( .A(n69), .ZN(n377) );
  INV_X1 U422 ( .A(n132), .ZN(n50) );
  NAND3_X1 U423 ( .A1(n50), .A2(n63), .A3(n141), .ZN(n387) );
  NAND3_X1 U424 ( .A1(n17), .A2(n231), .A3(n232), .ZN(n389) );
  INV_X1 U425 ( .A(n133), .ZN(n231) );
  NAND3_X1 U426 ( .A1(n401), .A2(n63), .A3(n141), .ZN(n400) );
  INV_X1 U427 ( .A(n103), .ZN(n141) );
  NAND2_X2 U428 ( .A1(A[21]), .A2(n409), .ZN(n88) );
  NAND2_X2 U429 ( .A1(A[17]), .A2(n410), .ZN(n91) );
  INV_X1 U430 ( .A(n94), .ZN(n392) );
endmodule


module ALU_N32 ( .FUNC({\FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] }), DATA1, 
        DATA2, OUTALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUTALU;
  input \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, \S[3] , net24446, net42480, net42491, net42492, net42493,
         net42498, net48162, net48160, net48158, net48196, net48194, net48192,
         net48190, net48188, net48186, net48200, net48198, net48204, net48202,
         net48208, net48206, net48212, net48210, net51555, net51683, net52829,
         net42478, net42477, net42476, net42426, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254;
  wire   [3:0] FUNC;
  wire   [31:0] Y_LOGIC;
  wire   [31:0] OUT_SHIFTER;
  wire   [31:0] L0;
  wire   [31:0] L1;
  wire   [31:0] L2;
  wire   [31:0] L3;

  BUF_X2 U5 ( .A(DATA2[15]), .Z(n69) );
  BUF_X1 U6 ( .A(DATA1[9]), .Z(n108) );
  INV_X1 U7 ( .A(n245), .ZN(n1) );
  CLKBUF_X3 U8 ( .A(DATA1[10]), .Z(n112) );
  CLKBUF_X3 U10 ( .A(DATA2[4]), .Z(n81) );
  INV_X1 U11 ( .A(n9), .ZN(n14) );
  BUF_X1 U12 ( .A(n40), .Z(net48204) );
  BUF_X1 U13 ( .A(n40), .Z(net48202) );
  AND2_X1 U14 ( .A1(Y_LOGIC[0]), .A2(net48206), .ZN(n2) );
  AND2_X1 U15 ( .A1(n35), .A2(n21), .ZN(n3) );
  INV_X1 U16 ( .A(n198), .ZN(n4) );
  BUF_X2 U17 ( .A(n89), .Z(n5) );
  AND2_X1 U18 ( .A1(n127), .A2(n130), .ZN(n6) );
  AND2_X1 U19 ( .A1(n175), .A2(n176), .ZN(n7) );
  OR2_X1 U20 ( .A1(n125), .A2(n8), .ZN(n9) );
  INV_X1 U21 ( .A(net51555), .ZN(n8) );
  AND2_X1 U22 ( .A1(N112), .A2(n14), .ZN(n124) );
  CLKBUF_X1 U23 ( .A(DATA2[25]), .Z(n15) );
  INV_X1 U24 ( .A(n242), .ZN(n16) );
  BUF_X1 U25 ( .A(DATA2[3]), .Z(n98) );
  CLKBUF_X1 U26 ( .A(DATA2[7]), .Z(n53) );
  INV_X1 U27 ( .A(DATA2[2]), .ZN(n17) );
  INV_X1 U28 ( .A(n17), .ZN(n18) );
  INV_X1 U29 ( .A(n196), .ZN(n19) );
  INV_X1 U30 ( .A(DATA1[3]), .ZN(n20) );
  CLKBUF_X1 U31 ( .A(FUNC[1]), .Z(n21) );
  CLKBUF_X3 U32 ( .A(DATA1[1]), .Z(n102) );
  BUF_X1 U33 ( .A(DATA1[20]), .Z(n22) );
  BUF_X2 U34 ( .A(DATA1[20]), .Z(n23) );
  NAND3_X1 U35 ( .A1(n174), .A2(n173), .A3(n7), .ZN(OUTALU[23]) );
  BUF_X1 U36 ( .A(DATA2[16]), .Z(n116) );
  NOR2_X1 U37 ( .A1(n24), .A2(n25), .ZN(n31) );
  AND2_X1 U38 ( .A1(N101), .A2(net48202), .ZN(n24) );
  NAND2_X1 U39 ( .A1(n32), .A2(n30), .ZN(n25) );
  INV_X1 U40 ( .A(net52829), .ZN(net42477) );
  CLKBUF_X1 U41 ( .A(DATA2[23]), .Z(n26) );
  CLKBUF_X1 U42 ( .A(DATA1[19]), .Z(n27) );
  BUF_X1 U43 ( .A(DATA1[19]), .Z(n28) );
  BUF_X2 U44 ( .A(DATA1[19]), .Z(n29) );
  NAND2_X1 U45 ( .A1(Y_LOGIC[22]), .A2(net48208), .ZN(n30) );
  NAND2_X1 U46 ( .A1(N69), .A2(net48200), .ZN(n32) );
  BUF_X1 U47 ( .A(DATA1[0]), .Z(n105) );
  AOI22_X1 U48 ( .A1(N62), .A2(n39), .B1(OUT_SHIFTER[15]), .B2(n34), .ZN(n160)
         );
  NAND2_X1 U49 ( .A1(n31), .A2(net42426), .ZN(OUTALU[22]) );
  NAND2_X1 U50 ( .A1(OUT_SHIFTER[22]), .A2(net48212), .ZN(net42426) );
  CLKBUF_X3 U51 ( .A(n34), .Z(net48212) );
  BUF_X2 U52 ( .A(n39), .Z(net48200) );
  BUF_X2 U53 ( .A(n33), .Z(net48208) );
  NAND2_X1 U54 ( .A1(net42476), .A2(net42477), .ZN(n34) );
  BUF_X2 U55 ( .A(n34), .Z(net48210) );
  NAND3_X1 U56 ( .A1(n21), .A2(net42478), .A3(n35), .ZN(net42476) );
  INV_X1 U57 ( .A(FUNC[0]), .ZN(n35) );
  AND3_X1 U58 ( .A1(net51683), .A2(n21), .A3(n35), .ZN(n40) );
  INV_X1 U59 ( .A(net42480), .ZN(net42478) );
  AND3_X1 U60 ( .A1(net51683), .A2(FUNC[0]), .A3(n36), .ZN(n39) );
  BUF_X2 U61 ( .A(n39), .Z(net48198) );
  INV_X1 U62 ( .A(FUNC[1]), .ZN(n36) );
  AND4_X2 U63 ( .A1(FUNC[3]), .A2(FUNC[0]), .A3(n36), .A4(net42498), .ZN(
        net52829) );
  AND2_X1 U64 ( .A1(N113), .A2(n36), .ZN(net42492) );
  NAND3_X1 U65 ( .A1(FUNC[2]), .A2(n36), .A3(net42491), .ZN(n37) );
  NAND2_X1 U66 ( .A1(n37), .A2(n38), .ZN(n33) );
  BUF_X2 U67 ( .A(n33), .Z(net48206) );
  NOR2_X1 U68 ( .A1(FUNC[0]), .A2(net42480), .ZN(net42493) );
  NAND2_X1 U69 ( .A1(net51555), .A2(net51683), .ZN(n38) );
  OAI21_X1 U70 ( .B1(FUNC[0]), .B2(n37), .A(n38), .ZN(\S[3] ) );
  INV_X1 U71 ( .A(n37), .ZN(net24446) );
  BUF_X1 U72 ( .A(DATA2[3]), .Z(n97) );
  CLKBUF_X1 U73 ( .A(DATA2[26]), .Z(n41) );
  CLKBUF_X1 U74 ( .A(DATA2[1]), .Z(n42) );
  CLKBUF_X1 U75 ( .A(DATA1[7]), .Z(n43) );
  BUF_X1 U76 ( .A(DATA1[25]), .Z(n59) );
  INV_X1 U77 ( .A(n200), .ZN(n44) );
  CLKBUF_X1 U78 ( .A(DATA2[21]), .Z(n45) );
  BUF_X2 U79 ( .A(DATA2[17]), .Z(n46) );
  CLKBUF_X1 U80 ( .A(DATA2[18]), .Z(n47) );
  INV_X1 U81 ( .A(n209), .ZN(n48) );
  BUF_X1 U82 ( .A(DATA1[22]), .Z(n49) );
  BUF_X1 U83 ( .A(DATA1[22]), .Z(n50) );
  BUF_X2 U84 ( .A(DATA1[22]), .Z(n51) );
  CLKBUF_X1 U85 ( .A(DATA1[4]), .Z(n52) );
  INV_X1 U86 ( .A(n118), .ZN(n54) );
  BUF_X1 U87 ( .A(DATA1[10]), .Z(n111) );
  CLKBUF_X1 U88 ( .A(DATA1[6]), .Z(n89) );
  CLKBUF_X1 U89 ( .A(DATA2[27]), .Z(n55) );
  CLKBUF_X1 U90 ( .A(DATA1[14]), .Z(n56) );
  CLKBUF_X1 U91 ( .A(DATA1[11]), .Z(n68) );
  CLKBUF_X3 U92 ( .A(DATA1[13]), .Z(n100) );
  CLKBUF_X1 U93 ( .A(DATA2[9]), .Z(n57) );
  INV_X1 U94 ( .A(n243), .ZN(n58) );
  BUF_X2 U95 ( .A(DATA1[25]), .Z(n60) );
  CLKBUF_X1 U96 ( .A(n57), .Z(n61) );
  BUF_X2 U97 ( .A(DATA1[0]), .Z(n106) );
  AND2_X1 U98 ( .A1(n77), .A2(n76), .ZN(n62) );
  AND2_X1 U99 ( .A1(n62), .A2(n75), .ZN(n186) );
  INV_X1 U100 ( .A(n214), .ZN(n63) );
  CLKBUF_X1 U101 ( .A(DATA1[5]), .Z(n64) );
  BUF_X1 U102 ( .A(DATA1[13]), .Z(n99) );
  INV_X1 U103 ( .A(n221), .ZN(n65) );
  INV_X1 U104 ( .A(n248), .ZN(n66) );
  INV_X1 U105 ( .A(n243), .ZN(n67) );
  INV_X1 U106 ( .A(n211), .ZN(n70) );
  INV_X1 U107 ( .A(n20), .ZN(n71) );
  INV_X1 U108 ( .A(n20), .ZN(n72) );
  INV_X1 U109 ( .A(n219), .ZN(n73) );
  CLKBUF_X1 U110 ( .A(DATA1[14]), .Z(n74) );
  NAND2_X1 U111 ( .A1(N106), .A2(net48202), .ZN(n75) );
  NAND2_X1 U112 ( .A1(Y_LOGIC[27]), .A2(net48208), .ZN(n76) );
  NAND2_X1 U113 ( .A1(N74), .A2(net48200), .ZN(n77) );
  BUF_X1 U114 ( .A(DATA2[4]), .Z(n80) );
  INV_X1 U115 ( .A(n222), .ZN(n78) );
  CLKBUF_X1 U116 ( .A(n97), .Z(n79) );
  INV_X1 U117 ( .A(n120), .ZN(n119) );
  INV_X1 U118 ( .A(n241), .ZN(n82) );
  NAND2_X1 U119 ( .A1(N108), .A2(net48202), .ZN(n83) );
  NAND2_X1 U120 ( .A1(Y_LOGIC[29]), .A2(net48208), .ZN(n84) );
  NAND2_X1 U121 ( .A1(N76), .A2(net48200), .ZN(n85) );
  AND3_X1 U122 ( .A1(n83), .A2(n84), .A3(n85), .ZN(n189) );
  NAND2_X1 U123 ( .A1(N78), .A2(net48198), .ZN(n86) );
  NAND2_X1 U124 ( .A1(N110), .A2(net48204), .ZN(n87) );
  NAND2_X1 U125 ( .A1(Y_LOGIC[31]), .A2(net48208), .ZN(n88) );
  AND3_X1 U126 ( .A1(n86), .A2(n87), .A3(n88), .ZN(n193) );
  NAND3_X1 U127 ( .A1(N111), .A2(n126), .A3(n3), .ZN(n127) );
  NAND3_X1 U128 ( .A1(n129), .A2(n128), .A3(n6), .ZN(OUTALU[0]) );
  NAND2_X1 U129 ( .A1(N77), .A2(net48198), .ZN(n90) );
  NAND2_X1 U130 ( .A1(N109), .A2(net48204), .ZN(n91) );
  NAND2_X1 U131 ( .A1(Y_LOGIC[30]), .A2(net48208), .ZN(n92) );
  AND3_X1 U132 ( .A1(n90), .A2(n91), .A3(n92), .ZN(n192) );
  NAND2_X1 U133 ( .A1(N75), .A2(net48198), .ZN(n93) );
  NAND2_X1 U134 ( .A1(N107), .A2(net48204), .ZN(n94) );
  NAND2_X1 U135 ( .A1(Y_LOGIC[28]), .A2(net48208), .ZN(n95) );
  AND3_X1 U136 ( .A1(n93), .A2(n94), .A3(n95), .ZN(n188) );
  CLKBUF_X1 U137 ( .A(DATA2[19]), .Z(n96) );
  NAND2_X1 U138 ( .A1(N73), .A2(net48198), .ZN(n181) );
  NAND2_X1 U139 ( .A1(N70), .A2(net48198), .ZN(n175) );
  NAND2_X1 U140 ( .A1(OUT_SHIFTER[0]), .A2(net48210), .ZN(n128) );
  NAND2_X1 U141 ( .A1(N105), .A2(net48202), .ZN(n184) );
  BUF_X2 U142 ( .A(net24446), .Z(net48190) );
  BUF_X2 U143 ( .A(net24446), .Z(net48188) );
  BUF_X2 U144 ( .A(net24446), .Z(net48194) );
  BUF_X2 U145 ( .A(net24446), .Z(net48192) );
  BUF_X2 U146 ( .A(net24446), .Z(net48186) );
  NAND2_X1 U147 ( .A1(N47), .A2(net48198), .ZN(n121) );
  NOR2_X1 U148 ( .A1(n124), .A2(n123), .ZN(n129) );
  NAND2_X1 U149 ( .A1(n122), .A2(n121), .ZN(n123) );
  NAND2_X1 U150 ( .A1(N79), .A2(net48202), .ZN(n122) );
  BUF_X2 U151 ( .A(\S[3] ), .Z(net48160) );
  BUF_X2 U152 ( .A(\S[3] ), .Z(net48158) );
  BUF_X2 U153 ( .A(\S[3] ), .Z(net48162) );
  AND2_X1 U154 ( .A1(net42491), .A2(net42498), .ZN(net51683) );
  INV_X1 U155 ( .A(n125), .ZN(n126) );
  NAND2_X1 U156 ( .A1(Y_LOGIC[23]), .A2(net48206), .ZN(n176) );
  NAND2_X1 U157 ( .A1(Y_LOGIC[26]), .A2(net48206), .ZN(n183) );
  AOI21_X1 U158 ( .B1(net42492), .B2(net42493), .A(n2), .ZN(n130) );
  AND2_X1 U159 ( .A1(FUNC[1]), .A2(FUNC[0]), .ZN(net51555) );
  CLKBUF_X1 U160 ( .A(DATA2[0]), .Z(n101) );
  BUF_X1 U161 ( .A(DATA2[28]), .Z(n103) );
  CLKBUF_X1 U162 ( .A(DATA2[28]), .Z(n104) );
  CLKBUF_X1 U163 ( .A(DATA1[0]), .Z(n107) );
  BUF_X2 U164 ( .A(DATA1[9]), .Z(n109) );
  BUF_X1 U165 ( .A(DATA1[9]), .Z(n110) );
  BUF_X2 U166 ( .A(DATA1[8]), .Z(n113) );
  BUF_X1 U167 ( .A(DATA1[8]), .Z(n114) );
  CLKBUF_X1 U168 ( .A(DATA2[30]), .Z(n115) );
  NAND2_X1 U169 ( .A1(OUT_SHIFTER[23]), .A2(net48210), .ZN(n174) );
  NAND4_X1 U170 ( .A1(n182), .A2(n183), .A3(n184), .A4(n181), .ZN(OUTALU[26])
         );
  NAND2_X1 U171 ( .A1(OUT_SHIFTER[26]), .A2(net48210), .ZN(n182) );
  NAND2_X1 U172 ( .A1(N102), .A2(net48202), .ZN(n173) );
  CLKBUF_X1 U173 ( .A(net24446), .Z(net48196) );
  INV_X1 U174 ( .A(n101), .ZN(n117) );
  INV_X1 U175 ( .A(DATA2[1]), .ZN(n118) );
  INV_X1 U176 ( .A(DATA2[2]), .ZN(n120) );
  INV_X1 U177 ( .A(FUNC[2]), .ZN(net42498) );
  INV_X1 U178 ( .A(FUNC[3]), .ZN(net42491) );
  INV_X1 U179 ( .A(DATA2[31]), .ZN(n225) );
  INV_X1 U180 ( .A(n115), .ZN(n226) );
  INV_X1 U181 ( .A(DATA2[29]), .ZN(n227) );
  INV_X1 U182 ( .A(n104), .ZN(n228) );
  INV_X1 U183 ( .A(DATA2[27]), .ZN(n229) );
  INV_X1 U184 ( .A(n41), .ZN(n230) );
  INV_X1 U185 ( .A(DATA2[25]), .ZN(n231) );
  INV_X1 U186 ( .A(DATA2[24]), .ZN(n232) );
  INV_X1 U187 ( .A(DATA2[23]), .ZN(n233) );
  INV_X1 U188 ( .A(DATA2[22]), .ZN(n234) );
  INV_X1 U189 ( .A(DATA2[21]), .ZN(n235) );
  INV_X1 U190 ( .A(DATA2[20]), .ZN(n236) );
  INV_X1 U191 ( .A(DATA2[19]), .ZN(n237) );
  INV_X1 U192 ( .A(n47), .ZN(n238) );
  INV_X1 U193 ( .A(n46), .ZN(n239) );
  INV_X1 U194 ( .A(DATA2[16]), .ZN(n240) );
  INV_X1 U195 ( .A(n69), .ZN(n241) );
  INV_X1 U196 ( .A(DATA2[14]), .ZN(n242) );
  INV_X1 U197 ( .A(DATA2[13]), .ZN(n243) );
  INV_X1 U198 ( .A(DATA2[12]), .ZN(n244) );
  INV_X1 U199 ( .A(DATA2[11]), .ZN(n245) );
  INV_X1 U200 ( .A(DATA2[10]), .ZN(n246) );
  INV_X1 U201 ( .A(n57), .ZN(n247) );
  INV_X1 U202 ( .A(DATA2[8]), .ZN(n248) );
  INV_X1 U203 ( .A(DATA2[7]), .ZN(n249) );
  INV_X1 U204 ( .A(DATA2[6]), .ZN(n250) );
  INV_X1 U205 ( .A(DATA2[5]), .ZN(n251) );
  INV_X1 U206 ( .A(n81), .ZN(n252) );
  INV_X1 U207 ( .A(n79), .ZN(n253) );
  INV_X1 U208 ( .A(DATA1[31]), .ZN(n195) );
  INV_X1 U209 ( .A(DATA1[30]), .ZN(n196) );
  INV_X1 U210 ( .A(DATA1[29]), .ZN(n197) );
  INV_X1 U211 ( .A(DATA1[28]), .ZN(n198) );
  INV_X1 U212 ( .A(DATA1[27]), .ZN(n199) );
  INV_X1 U213 ( .A(DATA1[26]), .ZN(n200) );
  INV_X1 U214 ( .A(n60), .ZN(n201) );
  INV_X1 U215 ( .A(DATA1[24]), .ZN(n202) );
  INV_X1 U216 ( .A(DATA1[23]), .ZN(n203) );
  INV_X1 U217 ( .A(n50), .ZN(n204) );
  INV_X1 U218 ( .A(DATA1[21]), .ZN(n205) );
  INV_X1 U219 ( .A(n22), .ZN(n206) );
  INV_X1 U220 ( .A(n28), .ZN(n207) );
  INV_X1 U221 ( .A(DATA1[18]), .ZN(n208) );
  INV_X1 U222 ( .A(DATA1[17]), .ZN(n209) );
  INV_X1 U223 ( .A(DATA1[16]), .ZN(n210) );
  INV_X1 U224 ( .A(DATA1[15]), .ZN(n211) );
  INV_X1 U225 ( .A(n74), .ZN(n212) );
  INV_X1 U226 ( .A(n100), .ZN(n213) );
  INV_X1 U227 ( .A(DATA1[12]), .ZN(n214) );
  INV_X1 U228 ( .A(n68), .ZN(n215) );
  INV_X1 U229 ( .A(n111), .ZN(n216) );
  INV_X1 U230 ( .A(n109), .ZN(n217) );
  INV_X1 U231 ( .A(n113), .ZN(n218) );
  INV_X1 U232 ( .A(n43), .ZN(n219) );
  INV_X1 U233 ( .A(n5), .ZN(n220) );
  INV_X1 U234 ( .A(n64), .ZN(n221) );
  INV_X1 U235 ( .A(DATA1[4]), .ZN(n222) );
  INV_X1 U236 ( .A(DATA1[2]), .ZN(n223) );
  INV_X1 U237 ( .A(n102), .ZN(n224) );
  INV_X1 U238 ( .A(n106), .ZN(n254) );
  NAND2_X1 U239 ( .A1(FUNC[3]), .A2(net42498), .ZN(net42480) );
  NAND2_X1 U240 ( .A1(FUNC[2]), .A2(net42491), .ZN(n125) );
  AOI22_X1 U241 ( .A1(OUT_SHIFTER[1]), .A2(net48210), .B1(N80), .B2(net48204), 
        .ZN(n132) );
  AOI22_X1 U242 ( .A1(Y_LOGIC[1]), .A2(net48206), .B1(N48), .B2(net48198), 
        .ZN(n131) );
  NAND2_X1 U243 ( .A1(n132), .A2(n131), .ZN(OUTALU[1]) );
  AOI22_X1 U244 ( .A1(OUT_SHIFTER[2]), .A2(net48212), .B1(N81), .B2(net48204), 
        .ZN(n134) );
  AOI22_X1 U245 ( .A1(Y_LOGIC[2]), .A2(net48206), .B1(N49), .B2(net48200), 
        .ZN(n133) );
  NAND2_X1 U246 ( .A1(n134), .A2(n133), .ZN(OUTALU[2]) );
  AOI22_X1 U247 ( .A1(OUT_SHIFTER[3]), .A2(net48212), .B1(N82), .B2(net48204), 
        .ZN(n136) );
  AOI22_X1 U248 ( .A1(Y_LOGIC[3]), .A2(net48206), .B1(N50), .B2(net48200), 
        .ZN(n135) );
  NAND2_X1 U249 ( .A1(n136), .A2(n135), .ZN(OUTALU[3]) );
  AOI22_X1 U250 ( .A1(OUT_SHIFTER[4]), .A2(net48212), .B1(N83), .B2(net48204), 
        .ZN(n138) );
  AOI22_X1 U251 ( .A1(Y_LOGIC[4]), .A2(net48206), .B1(N51), .B2(net48200), 
        .ZN(n137) );
  NAND2_X1 U252 ( .A1(n138), .A2(n137), .ZN(OUTALU[4]) );
  AOI22_X1 U253 ( .A1(OUT_SHIFTER[5]), .A2(net48212), .B1(N84), .B2(net48204), 
        .ZN(n140) );
  AOI22_X1 U254 ( .A1(Y_LOGIC[5]), .A2(net48206), .B1(N52), .B2(net48200), 
        .ZN(n139) );
  NAND2_X1 U255 ( .A1(n140), .A2(n139), .ZN(OUTALU[5]) );
  AOI22_X1 U256 ( .A1(OUT_SHIFTER[6]), .A2(net48210), .B1(N85), .B2(net48204), 
        .ZN(n142) );
  AOI22_X1 U257 ( .A1(Y_LOGIC[6]), .A2(net48206), .B1(N53), .B2(net48200), 
        .ZN(n141) );
  NAND2_X1 U258 ( .A1(n142), .A2(n141), .ZN(OUTALU[6]) );
  AOI22_X1 U259 ( .A1(OUT_SHIFTER[7]), .A2(net48212), .B1(N86), .B2(net48204), 
        .ZN(n144) );
  AOI22_X1 U260 ( .A1(Y_LOGIC[7]), .A2(net48206), .B1(N54), .B2(net48200), 
        .ZN(n143) );
  NAND2_X1 U261 ( .A1(n144), .A2(n143), .ZN(OUTALU[7]) );
  AOI22_X1 U262 ( .A1(OUT_SHIFTER[8]), .A2(net48210), .B1(N87), .B2(net48202), 
        .ZN(n146) );
  AOI22_X1 U263 ( .A1(Y_LOGIC[8]), .A2(net48206), .B1(N55), .B2(net48198), 
        .ZN(n145) );
  NAND2_X1 U264 ( .A1(n146), .A2(n145), .ZN(OUTALU[8]) );
  AOI22_X1 U265 ( .A1(OUT_SHIFTER[9]), .A2(net48212), .B1(N88), .B2(net48202), 
        .ZN(n148) );
  AOI22_X1 U266 ( .A1(Y_LOGIC[9]), .A2(net48206), .B1(N56), .B2(net48200), 
        .ZN(n147) );
  NAND2_X1 U267 ( .A1(n148), .A2(n147), .ZN(OUTALU[9]) );
  AOI22_X1 U268 ( .A1(OUT_SHIFTER[10]), .A2(net48212), .B1(N89), .B2(net48202), 
        .ZN(n150) );
  AOI22_X1 U269 ( .A1(Y_LOGIC[10]), .A2(net48206), .B1(N57), .B2(net48200), 
        .ZN(n149) );
  NAND2_X1 U270 ( .A1(n150), .A2(n149), .ZN(OUTALU[10]) );
  AOI22_X1 U271 ( .A1(OUT_SHIFTER[11]), .A2(net48210), .B1(N90), .B2(net48202), 
        .ZN(n152) );
  AOI22_X1 U272 ( .A1(Y_LOGIC[11]), .A2(net48206), .B1(N58), .B2(net48200), 
        .ZN(n151) );
  NAND2_X1 U273 ( .A1(n152), .A2(n151), .ZN(OUTALU[11]) );
  AOI22_X1 U274 ( .A1(OUT_SHIFTER[12]), .A2(net48210), .B1(N91), .B2(net48202), 
        .ZN(n154) );
  AOI22_X1 U275 ( .A1(Y_LOGIC[12]), .A2(net48206), .B1(N59), .B2(net48200), 
        .ZN(n153) );
  NAND2_X1 U276 ( .A1(n154), .A2(n153), .ZN(OUTALU[12]) );
  AOI22_X1 U277 ( .A1(OUT_SHIFTER[13]), .A2(net48210), .B1(N92), .B2(net48202), 
        .ZN(n156) );
  AOI22_X1 U278 ( .A1(Y_LOGIC[13]), .A2(net48208), .B1(N60), .B2(net48198), 
        .ZN(n155) );
  NAND2_X1 U279 ( .A1(n156), .A2(n155), .ZN(OUTALU[13]) );
  AOI22_X1 U280 ( .A1(OUT_SHIFTER[14]), .A2(net48210), .B1(N93), .B2(net48202), 
        .ZN(n158) );
  AOI22_X1 U281 ( .A1(Y_LOGIC[14]), .A2(net48206), .B1(N61), .B2(net48198), 
        .ZN(n157) );
  NAND2_X1 U282 ( .A1(n158), .A2(n157), .ZN(OUTALU[14]) );
  AOI22_X1 U283 ( .A1(N94), .A2(net48202), .B1(Y_LOGIC[15]), .B2(net48208), 
        .ZN(n159) );
  NAND2_X1 U284 ( .A1(n160), .A2(n159), .ZN(OUTALU[15]) );
  AOI22_X1 U285 ( .A1(OUT_SHIFTER[16]), .A2(net48210), .B1(N95), .B2(net48202), 
        .ZN(n162) );
  AOI22_X1 U286 ( .A1(Y_LOGIC[16]), .A2(net48206), .B1(N63), .B2(net48198), 
        .ZN(n161) );
  NAND2_X1 U287 ( .A1(n162), .A2(n161), .ZN(OUTALU[16]) );
  AOI22_X1 U288 ( .A1(OUT_SHIFTER[17]), .A2(net48210), .B1(N96), .B2(net48202), 
        .ZN(n164) );
  AOI22_X1 U289 ( .A1(Y_LOGIC[17]), .A2(net48206), .B1(N64), .B2(net48198), 
        .ZN(n163) );
  NAND2_X1 U290 ( .A1(n164), .A2(n163), .ZN(OUTALU[17]) );
  AOI22_X1 U291 ( .A1(OUT_SHIFTER[18]), .A2(net48210), .B1(N97), .B2(net48204), 
        .ZN(n166) );
  AOI22_X1 U292 ( .A1(Y_LOGIC[18]), .A2(net48208), .B1(N65), .B2(net48198), 
        .ZN(n165) );
  NAND2_X1 U293 ( .A1(n166), .A2(n165), .ZN(OUTALU[18]) );
  AOI222_X1 U294 ( .A1(OUT_SHIFTER[19]), .A2(net48210), .B1(Y_LOGIC[19]), .B2(
        net48208), .C1(N66), .C2(net48200), .ZN(n168) );
  NAND2_X1 U295 ( .A1(N98), .A2(net48202), .ZN(n167) );
  NAND2_X1 U296 ( .A1(n167), .A2(n168), .ZN(OUTALU[19]) );
  AOI22_X1 U297 ( .A1(OUT_SHIFTER[20]), .A2(net48210), .B1(N99), .B2(net48204), 
        .ZN(n170) );
  AOI22_X1 U298 ( .A1(Y_LOGIC[20]), .A2(net48208), .B1(N67), .B2(net48198), 
        .ZN(n169) );
  NAND2_X1 U299 ( .A1(n170), .A2(n169), .ZN(OUTALU[20]) );
  AOI22_X1 U300 ( .A1(OUT_SHIFTER[21]), .A2(net48210), .B1(N100), .B2(net48204), .ZN(n172) );
  AOI22_X1 U301 ( .A1(Y_LOGIC[21]), .A2(net48208), .B1(N68), .B2(net48198), 
        .ZN(n171) );
  NAND2_X1 U302 ( .A1(n172), .A2(n171), .ZN(OUTALU[21]) );
  AOI22_X1 U303 ( .A1(OUT_SHIFTER[24]), .A2(net48210), .B1(N71), .B2(net48198), 
        .ZN(n178) );
  AOI22_X1 U304 ( .A1(N103), .A2(net48202), .B1(Y_LOGIC[24]), .B2(net48208), 
        .ZN(n177) );
  NAND2_X1 U305 ( .A1(n178), .A2(n177), .ZN(OUTALU[24]) );
  AOI22_X1 U306 ( .A1(OUT_SHIFTER[25]), .A2(net48210), .B1(N104), .B2(net48204), .ZN(n180) );
  AOI22_X1 U307 ( .A1(Y_LOGIC[25]), .A2(net48208), .B1(N72), .B2(net48198), 
        .ZN(n179) );
  NAND2_X1 U308 ( .A1(n180), .A2(n179), .ZN(OUTALU[25]) );
  NAND2_X1 U309 ( .A1(OUT_SHIFTER[27]), .A2(net48212), .ZN(n185) );
  NAND2_X1 U310 ( .A1(n185), .A2(n186), .ZN(OUTALU[27]) );
  NAND2_X1 U311 ( .A1(OUT_SHIFTER[28]), .A2(net48212), .ZN(n187) );
  NAND2_X1 U312 ( .A1(n187), .A2(n188), .ZN(OUTALU[28]) );
  NAND2_X1 U313 ( .A1(OUT_SHIFTER[29]), .A2(net48212), .ZN(n190) );
  NAND2_X1 U314 ( .A1(n190), .A2(n189), .ZN(OUTALU[29]) );
  NAND2_X1 U315 ( .A1(OUT_SHIFTER[30]), .A2(net48212), .ZN(n191) );
  NAND2_X1 U316 ( .A1(n192), .A2(n191), .ZN(OUTALU[30]) );
  NAND2_X1 U317 ( .A1(OUT_SHIFTER[31]), .A2(net48212), .ZN(n194) );
  NAND2_X1 U318 ( .A1(n193), .A2(n194), .ZN(OUTALU[31]) );
  NAND3_0 NAND31I_1 ( .A(n254), .B(n117), .C(1'b0), .Y(L0[0]) );
  NAND3_127 NAND31I_2 ( .A(n224), .B(n118), .C(1'b0), .Y(L0[1]) );
  NAND3_126 NAND31I_3 ( .A(n223), .B(n120), .C(1'b0), .Y(L0[2]) );
  NAND3_125 NAND31I_4 ( .A(n20), .B(n253), .C(1'b0), .Y(L0[3]) );
  NAND3_124 NAND31I_5 ( .A(n222), .B(n252), .C(1'b0), .Y(L0[4]) );
  NAND3_123 NAND31I_6 ( .A(n221), .B(n251), .C(1'b0), .Y(L0[5]) );
  NAND3_122 NAND31I_7 ( .A(n220), .B(n250), .C(1'b0), .Y(L0[6]) );
  NAND3_121 NAND31I_8 ( .A(n219), .B(n249), .C(1'b0), .Y(L0[7]) );
  NAND3_120 NAND31I_9 ( .A(n218), .B(n248), .C(1'b0), .Y(L0[8]) );
  NAND3_119 NAND31I_10 ( .A(n217), .B(n247), .C(1'b0), .Y(L0[9]) );
  NAND3_118 NAND31I_11 ( .A(n216), .B(n246), .C(1'b0), .Y(L0[10]) );
  NAND3_117 NAND31I_12 ( .A(n215), .B(n245), .C(1'b0), .Y(L0[11]) );
  NAND3_116 NAND31I_13 ( .A(n214), .B(n244), .C(1'b0), .Y(L0[12]) );
  NAND3_115 NAND31I_14 ( .A(n213), .B(n243), .C(1'b0), .Y(L0[13]) );
  NAND3_114 NAND31I_15 ( .A(n212), .B(n242), .C(1'b0), .Y(L0[14]) );
  NAND3_113 NAND31I_16 ( .A(n211), .B(n241), .C(1'b0), .Y(L0[15]) );
  NAND3_112 NAND31I_17 ( .A(n210), .B(n240), .C(1'b0), .Y(L0[16]) );
  NAND3_111 NAND31I_18 ( .A(n209), .B(n239), .C(1'b0), .Y(L0[17]) );
  NAND3_110 NAND31I_19 ( .A(n208), .B(n238), .C(1'b0), .Y(L0[18]) );
  NAND3_109 NAND31I_20 ( .A(n207), .B(n237), .C(1'b0), .Y(L0[19]) );
  NAND3_108 NAND31I_21 ( .A(n206), .B(n236), .C(1'b0), .Y(L0[20]) );
  NAND3_107 NAND31I_22 ( .A(n205), .B(n235), .C(1'b0), .Y(L0[21]) );
  NAND3_106 NAND31I_23 ( .A(n204), .B(n234), .C(1'b0), .Y(L0[22]) );
  NAND3_105 NAND31I_24 ( .A(n203), .B(n233), .C(1'b0), .Y(L0[23]) );
  NAND3_104 NAND31I_25 ( .A(n202), .B(n232), .C(1'b0), .Y(L0[24]) );
  NAND3_103 NAND31I_26 ( .A(n201), .B(n231), .C(1'b0), .Y(L0[25]) );
  NAND3_102 NAND31I_27 ( .A(n200), .B(n230), .C(1'b0), .Y(L0[26]) );
  NAND3_101 NAND31I_28 ( .A(n199), .B(n229), .C(1'b0), .Y(L0[27]) );
  NAND3_100 NAND31I_29 ( .A(n198), .B(n228), .C(1'b0), .Y(L0[28]) );
  NAND3_99 NAND31I_30 ( .A(n197), .B(n227), .C(1'b0), .Y(L0[29]) );
  NAND3_98 NAND31I_31 ( .A(n196), .B(n226), .C(1'b0), .Y(L0[30]) );
  NAND3_97 NAND31I_32 ( .A(n195), .B(n225), .C(1'b0), .Y(L0[31]) );
  NAND3_96 NAND31I_1_0 ( .A(n254), .B(n101), .C(net48186), .Y(L1[0]) );
  NAND3_95 NAND31I_2_0 ( .A(n224), .B(n54), .C(net48186), .Y(L1[1]) );
  NAND3_94 NAND31I_3_0 ( .A(n223), .B(n119), .C(net48186), .Y(L1[2]) );
  NAND3_93 NAND31I_4_0 ( .A(n20), .B(n79), .C(net48186), .Y(L1[3]) );
  NAND3_92 NAND31I_5_0 ( .A(n222), .B(n81), .C(net48186), .Y(L1[4]) );
  NAND3_91 NAND31I_6_0 ( .A(n221), .B(DATA2[5]), .C(net48186), .Y(L1[5]) );
  NAND3_90 NAND31I_7_0 ( .A(n220), .B(DATA2[6]), .C(net48186), .Y(L1[6]) );
  NAND3_89 NAND31I_8_0 ( .A(n219), .B(DATA2[7]), .C(net48186), .Y(L1[7]) );
  NAND3_88 NAND31I_9_0 ( .A(n218), .B(n66), .C(net48186), .Y(L1[8]) );
  NAND3_87 NAND31I_10_0 ( .A(n217), .B(n61), .C(net48186), .Y(L1[9]) );
  NAND3_86 NAND31I_11_0 ( .A(n216), .B(DATA2[10]), .C(net48186), .Y(L1[10]) );
  NAND3_85 NAND31I_12_0 ( .A(n215), .B(n1), .C(net48186), .Y(L1[11]) );
  NAND3_84 NAND31I_13_0 ( .A(n214), .B(DATA2[12]), .C(net48188), .Y(L1[12]) );
  NAND3_83 NAND31I_14_0 ( .A(n213), .B(n67), .C(net48188), .Y(L1[13]) );
  NAND3_82 NAND31I_15_0 ( .A(n212), .B(n16), .C(net48188), .Y(L1[14]) );
  NAND3_81 NAND31I_16_0 ( .A(n211), .B(n82), .C(net48188), .Y(L1[15]) );
  NAND3_80 NAND31I_17_0 ( .A(n210), .B(DATA2[16]), .C(net48188), .Y(L1[16]) );
  NAND3_79 NAND31I_18_0 ( .A(n209), .B(n46), .C(net48188), .Y(L1[17]) );
  NAND3_78 NAND31I_19_0 ( .A(n208), .B(n47), .C(net48188), .Y(L1[18]) );
  NAND3_77 NAND31I_20_0 ( .A(n207), .B(n96), .C(net48188), .Y(L1[19]) );
  NAND3_76 NAND31I_21_0 ( .A(n206), .B(DATA2[20]), .C(net48188), .Y(L1[20]) );
  NAND3_75 NAND31I_22_0 ( .A(n205), .B(DATA2[21]), .C(net48188), .Y(L1[21]) );
  NAND3_74 NAND31I_23_0 ( .A(n204), .B(DATA2[22]), .C(net48188), .Y(L1[22]) );
  NAND3_73 NAND31I_24_0 ( .A(n203), .B(DATA2[23]), .C(net48188), .Y(L1[23]) );
  NAND3_72 NAND31I_25_0 ( .A(n202), .B(DATA2[24]), .C(net48190), .Y(L1[24]) );
  NAND3_71 NAND31I_26_0 ( .A(n201), .B(n15), .C(net48190), .Y(L1[25]) );
  NAND3_70 NAND31I_27_0 ( .A(n200), .B(n41), .C(net48190), .Y(L1[26]) );
  NAND3_69 NAND31I_28_0 ( .A(n199), .B(DATA2[27]), .C(net48190), .Y(L1[27]) );
  NAND3_68 NAND31I_29_0 ( .A(n198), .B(n104), .C(net48190), .Y(L1[28]) );
  NAND3_67 NAND31I_30_0 ( .A(n197), .B(DATA2[29]), .C(net48190), .Y(L1[29]) );
  NAND3_66 NAND31I_31_0 ( .A(n196), .B(n115), .C(net48190), .Y(L1[30]) );
  NAND3_65 NAND31I_32_0 ( .A(n195), .B(DATA2[31]), .C(net48190), .Y(L1[31]) );
  NAND3_64 NAND31I_1_1 ( .A(n107), .B(n117), .C(net48190), .Y(L2[0]) );
  NAND3_63 NAND31I_2_1 ( .A(n102), .B(n118), .C(net48190), .Y(L2[1]) );
  NAND3_62 NAND31I_3_1 ( .A(DATA1[2]), .B(n120), .C(net48190), .Y(L2[2]) );
  NAND3_61 NAND31I_4_1 ( .A(n72), .B(n253), .C(net48190), .Y(L2[3]) );
  NAND3_60 NAND31I_5_1 ( .A(n78), .B(n252), .C(net48192), .Y(L2[4]) );
  NAND3_59 NAND31I_6_1 ( .A(n64), .B(n251), .C(net48192), .Y(L2[5]) );
  NAND3_58 NAND31I_7_1 ( .A(n5), .B(n250), .C(net48192), .Y(L2[6]) );
  NAND3_57 NAND31I_8_1 ( .A(n73), .B(n249), .C(net48192), .Y(L2[7]) );
  NAND3_56 NAND31I_9_1 ( .A(n114), .B(n248), .C(net48192), .Y(L2[8]) );
  NAND3_55 NAND31I_10_1 ( .A(n110), .B(n247), .C(net48192), .Y(L2[9]) );
  NAND3_54 NAND31I_11_1 ( .A(n112), .B(n246), .C(net48192), .Y(L2[10]) );
  NAND3_53 NAND31I_12_1 ( .A(n68), .B(n245), .C(net48192), .Y(L2[11]) );
  NAND3_52 NAND31I_13_1 ( .A(n63), .B(n244), .C(net48192), .Y(L2[12]) );
  NAND3_51 NAND31I_14_1 ( .A(n100), .B(n243), .C(net48192), .Y(L2[13]) );
  NAND3_50 NAND31I_15_1 ( .A(n74), .B(n242), .C(net48192), .Y(L2[14]) );
  NAND3_49 NAND31I_16_1 ( .A(n70), .B(n241), .C(net48192), .Y(L2[15]) );
  NAND3_48 NAND31I_17_1 ( .A(DATA1[16]), .B(n240), .C(net48194), .Y(L2[16]) );
  NAND3_47 NAND31I_18_1 ( .A(n48), .B(n239), .C(net48194), .Y(L2[17]) );
  NAND3_46 NAND31I_19_1 ( .A(DATA1[18]), .B(n238), .C(net48194), .Y(L2[18]) );
  NAND3_45 NAND31I_20_1 ( .A(n29), .B(n237), .C(net48194), .Y(L2[19]) );
  NAND3_44 NAND31I_21_1 ( .A(n23), .B(n236), .C(net48194), .Y(L2[20]) );
  NAND3_43 NAND31I_22_1 ( .A(DATA1[21]), .B(n235), .C(net48194), .Y(L2[21]) );
  NAND3_42 NAND31I_23_1 ( .A(n51), .B(n234), .C(net48194), .Y(L2[22]) );
  NAND3_41 NAND31I_24_1 ( .A(DATA1[23]), .B(n233), .C(net48194), .Y(L2[23]) );
  NAND3_40 NAND31I_25_1 ( .A(DATA1[24]), .B(n232), .C(net48194), .Y(L2[24]) );
  NAND3_39 NAND31I_26_1 ( .A(n60), .B(n231), .C(net48194), .Y(L2[25]) );
  NAND3_38 NAND31I_27_1 ( .A(n44), .B(n230), .C(net48194), .Y(L2[26]) );
  NAND3_37 NAND31I_28_1 ( .A(DATA1[27]), .B(n229), .C(net48194), .Y(L2[27]) );
  NAND3_36 NAND31I_29_1 ( .A(n4), .B(n228), .C(net48196), .Y(L2[28]) );
  NAND3_35 NAND31I_30_1 ( .A(DATA1[29]), .B(n227), .C(net48196), .Y(L2[29]) );
  NAND3_34 NAND31I_31_1 ( .A(n19), .B(n226), .C(net48196), .Y(L2[30]) );
  NAND3_33 NAND31I_32_1 ( .A(DATA1[31]), .B(n225), .C(net48196), .Y(L2[31]) );
  NAND3_32 NAND31I_1_2 ( .A(n106), .B(n101), .C(net48158), .Y(L3[0]) );
  NAND3_31 NAND31I_2_2 ( .A(n102), .B(n54), .C(net48158), .Y(L3[1]) );
  NAND3_30 NAND31I_3_2 ( .A(DATA1[2]), .B(n119), .C(net48158), .Y(L3[2]) );
  NAND3_29 NAND31I_4_2 ( .A(n72), .B(n79), .C(net48158), .Y(L3[3]) );
  NAND3_28 NAND31I_5_2 ( .A(n78), .B(n81), .C(net48158), .Y(L3[4]) );
  NAND3_27 NAND31I_6_2 ( .A(n64), .B(DATA2[5]), .C(net48158), .Y(L3[5]) );
  NAND3_26 NAND31I_7_2 ( .A(n5), .B(DATA2[6]), .C(net48158), .Y(L3[6]) );
  NAND3_25 NAND31I_8_2 ( .A(n73), .B(n53), .C(net48158), .Y(L3[7]) );
  NAND3_24 NAND31I_9_2 ( .A(n113), .B(n66), .C(net48158), .Y(L3[8]) );
  NAND3_23 NAND31I_10_2 ( .A(n109), .B(n61), .C(net48158), .Y(L3[9]) );
  NAND3_22 NAND31I_11_2 ( .A(n111), .B(DATA2[10]), .C(net48158), .Y(L3[10]) );
  NAND3_21 NAND31I_12_2 ( .A(n68), .B(n1), .C(net48158), .Y(L3[11]) );
  NAND3_20 NAND31I_13_2 ( .A(n63), .B(DATA2[12]), .C(net48160), .Y(L3[12]) );
  NAND3_19 NAND31I_14_2 ( .A(n100), .B(n67), .C(net48160), .Y(L3[13]) );
  NAND3_18 NAND31I_15_2 ( .A(n56), .B(n16), .C(net48160), .Y(L3[14]) );
  NAND3_17 NAND31I_16_2 ( .A(n70), .B(n82), .C(net48160), .Y(L3[15]) );
  NAND3_16 NAND31I_17_2 ( .A(DATA1[16]), .B(n116), .C(net48160), .Y(L3[16]) );
  NAND3_15 NAND31I_18_2 ( .A(n48), .B(n46), .C(net48160), .Y(L3[17]) );
  NAND3_14 NAND31I_19_2 ( .A(DATA1[18]), .B(n47), .C(net48160), .Y(L3[18]) );
  NAND3_13 NAND31I_20_2 ( .A(n28), .B(DATA2[19]), .C(net48160), .Y(L3[19]) );
  NAND3_12 NAND31I_21_2 ( .A(n22), .B(DATA2[20]), .C(net48160), .Y(L3[20]) );
  NAND3_11 NAND31I_22_2 ( .A(DATA1[21]), .B(DATA2[21]), .C(net48160), .Y(
        L3[21]) );
  NAND3_10 NAND31I_23_2 ( .A(n50), .B(DATA2[22]), .C(net48160), .Y(L3[22]) );
  NAND3_9 NAND31I_24_2 ( .A(DATA1[23]), .B(DATA2[23]), .C(net48160), .Y(L3[23]) );
  NAND3_8 NAND31I_25_2 ( .A(DATA1[24]), .B(DATA2[24]), .C(net48162), .Y(L3[24]) );
  NAND3_7 NAND31I_26_2 ( .A(n60), .B(n15), .C(net48162), .Y(L3[25]) );
  NAND3_6 NAND31I_27_2 ( .A(n44), .B(n41), .C(net48162), .Y(L3[26]) );
  NAND3_5 NAND31I_28_2 ( .A(DATA1[27]), .B(DATA2[27]), .C(net48162), .Y(L3[27]) );
  NAND3_4 NAND31I_29_2 ( .A(n4), .B(n104), .C(net48162), .Y(L3[28]) );
  NAND3_3 NAND31I_30_2 ( .A(DATA1[29]), .B(DATA2[29]), .C(net48162), .Y(L3[29]) );
  NAND3_2 NAND31I_31_2 ( .A(n19), .B(n115), .C(net48162), .Y(L3[30]) );
  NAND3_1 NAND31I_32_2 ( .A(DATA1[31]), .B(DATA2[31]), .C(net48162), .Y(L3[31]) );
  NAND4_0 NAND41I_1 ( .A(L0[0]), .B(L1[0]), .C(L2[0]), .D(L3[0]), .Y(
        Y_LOGIC[0]) );
  NAND4_31 NAND41I_2 ( .A(L0[1]), .B(L1[1]), .C(L2[1]), .D(L3[1]), .Y(
        Y_LOGIC[1]) );
  NAND4_30 NAND41I_3 ( .A(L0[2]), .B(L1[2]), .C(L2[2]), .D(L3[2]), .Y(
        Y_LOGIC[2]) );
  NAND4_29 NAND41I_4 ( .A(L0[3]), .B(L1[3]), .C(L2[3]), .D(L3[3]), .Y(
        Y_LOGIC[3]) );
  NAND4_28 NAND41I_5 ( .A(L0[4]), .B(L1[4]), .C(L2[4]), .D(L3[4]), .Y(
        Y_LOGIC[4]) );
  NAND4_27 NAND41I_6 ( .A(L0[5]), .B(L1[5]), .C(L2[5]), .D(L3[5]), .Y(
        Y_LOGIC[5]) );
  NAND4_26 NAND41I_7 ( .A(L0[6]), .B(L1[6]), .C(L2[6]), .D(L3[6]), .Y(
        Y_LOGIC[6]) );
  NAND4_25 NAND41I_8 ( .A(L0[7]), .B(L1[7]), .C(L2[7]), .D(L3[7]), .Y(
        Y_LOGIC[7]) );
  NAND4_24 NAND41I_9 ( .A(L0[8]), .B(L1[8]), .C(L2[8]), .D(L3[8]), .Y(
        Y_LOGIC[8]) );
  NAND4_23 NAND41I_10 ( .A(L0[9]), .B(L1[9]), .C(L2[9]), .D(L3[9]), .Y(
        Y_LOGIC[9]) );
  NAND4_22 NAND41I_11 ( .A(L0[10]), .B(L1[10]), .C(L2[10]), .D(L3[10]), .Y(
        Y_LOGIC[10]) );
  NAND4_21 NAND41I_12 ( .A(L0[11]), .B(L1[11]), .C(L2[11]), .D(L3[11]), .Y(
        Y_LOGIC[11]) );
  NAND4_20 NAND41I_13 ( .A(L0[12]), .B(L1[12]), .C(L2[12]), .D(L3[12]), .Y(
        Y_LOGIC[12]) );
  NAND4_19 NAND41I_14 ( .A(L0[13]), .B(L1[13]), .C(L2[13]), .D(L3[13]), .Y(
        Y_LOGIC[13]) );
  NAND4_18 NAND41I_15 ( .A(L0[14]), .B(L1[14]), .C(L2[14]), .D(L3[14]), .Y(
        Y_LOGIC[14]) );
  NAND4_17 NAND41I_16 ( .A(L0[15]), .B(L1[15]), .C(L2[15]), .D(L3[15]), .Y(
        Y_LOGIC[15]) );
  NAND4_16 NAND41I_17 ( .A(L0[16]), .B(L1[16]), .C(L2[16]), .D(L3[16]), .Y(
        Y_LOGIC[16]) );
  NAND4_15 NAND41I_18 ( .A(L0[17]), .B(L1[17]), .C(L2[17]), .D(L3[17]), .Y(
        Y_LOGIC[17]) );
  NAND4_14 NAND41I_19 ( .A(L0[18]), .B(L1[18]), .C(L2[18]), .D(L3[18]), .Y(
        Y_LOGIC[18]) );
  NAND4_13 NAND41I_20 ( .A(L0[19]), .B(L1[19]), .C(L2[19]), .D(L3[19]), .Y(
        Y_LOGIC[19]) );
  NAND4_12 NAND41I_21 ( .A(L0[20]), .B(L1[20]), .C(L2[20]), .D(L3[20]), .Y(
        Y_LOGIC[20]) );
  NAND4_11 NAND41I_22 ( .A(L0[21]), .B(L1[21]), .C(L2[21]), .D(L3[21]), .Y(
        Y_LOGIC[21]) );
  NAND4_10 NAND41I_23 ( .A(L0[22]), .B(L1[22]), .C(L2[22]), .D(L3[22]), .Y(
        Y_LOGIC[22]) );
  NAND4_9 NAND41I_24 ( .A(L0[23]), .B(L1[23]), .C(L2[23]), .D(L3[23]), .Y(
        Y_LOGIC[23]) );
  NAND4_8 NAND41I_25 ( .A(L0[24]), .B(L1[24]), .C(L2[24]), .D(L3[24]), .Y(
        Y_LOGIC[24]) );
  NAND4_7 NAND41I_26 ( .A(L0[25]), .B(L1[25]), .C(L2[25]), .D(L3[25]), .Y(
        Y_LOGIC[25]) );
  NAND4_6 NAND41I_27 ( .A(L0[26]), .B(L1[26]), .C(L2[26]), .D(L3[26]), .Y(
        Y_LOGIC[26]) );
  NAND4_5 NAND41I_28 ( .A(L0[27]), .B(L1[27]), .C(L2[27]), .D(L3[27]), .Y(
        Y_LOGIC[27]) );
  NAND4_4 NAND41I_29 ( .A(L0[28]), .B(L1[28]), .C(L2[28]), .D(L3[28]), .Y(
        Y_LOGIC[28]) );
  NAND4_3 NAND41I_30 ( .A(L0[29]), .B(L1[29]), .C(L2[29]), .D(L3[29]), .Y(
        Y_LOGIC[29]) );
  NAND4_2 NAND41I_31 ( .A(L0[30]), .B(L1[30]), .C(L2[30]), .D(L3[30]), .Y(
        Y_LOGIC[30]) );
  NAND4_1 NAND41I_32 ( .A(L0[31]), .B(L1[31]), .C(L2[31]), .D(L3[31]), .Y(
        Y_LOGIC[31]) );
  BARREL_SHIFTER_N32 SHIFTER ( .CONF(net52829), .DATA1({DATA1[31:26], n60, 
        DATA1[24:23], n50, DATA1[21], n22, n28, DATA1[18], n48, DATA1[16:15], 
        n74, n100, DATA1[12], n68, n112, n109, n113, n43, n5, n64, n52, n71, 
        DATA1[2], n102, n106}), .DATA2({DATA2[31], n115, DATA2[29], n104, 
        DATA2[27], n41, n15, DATA2[24], n26, DATA2[22], n45, DATA2[20], n96, 
        n47, n46, DATA2[16], n82, n16, n67, DATA2[12], n1, DATA2[10], n61, n66, 
        DATA2[7:5], n80, n98, n18, n42, n101}), .OUTPUT(OUT_SHIFTER) );
  ALU_N32_DW01_sub_2 sub_66 ( .A({DATA1[31:26], n60, DATA1[24:23], n51, 
        DATA1[21], n23, n27, DATA1[18:10], n108, n113, DATA1[7:1], n105}), .B(
        {DATA2[31], n115, DATA2[29], n104, DATA2[27:18], n46, DATA2[16], n69, 
        DATA2[14:5], n81, n97, DATA2[2:0]}), .CI(1'b0), .DIFF({N110, N109, 
        N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, 
        N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, 
        N82, N81, N80, N79}) );
  ALU_N32_DW01_cmp6_4 ne_72 ( .A({DATA1[31], n19, DATA1[29], n4, DATA1[27], 
        n44, n60, DATA1[24:23], n51, DATA1[21], n23, n29, DATA1[18], n48, 
        DATA1[16], n70, n74, n100, n63, n68, n112, n110, n114, n73, n5, n65, 
        n78, n72, DATA1[2], n102, n107}), .B({DATA2[31], n115, DATA2[29], n104, 
        n55, n41, n15, DATA2[24:19], n47, n46, n116, n82, n16, n67, DATA2[12], 
        n1, DATA2[10], n57, n66, n53, DATA2[6:5], n81, n79, n119, n54, n101}), 
        .TC(1'b0), .NE(N113) );
  ALU_N32_DW01_add_4 add_65 ( .A({DATA1[31:26], n59, DATA1[24:23], n51, 
        DATA1[21], n23, n29, DATA1[18:14], n99, DATA1[12:11], n111, n109, 
        DATA1[8:1], n106}), .B({DATA2[31], n115, DATA2[29], n104, DATA2[27:5], 
        n81, n97, DATA2[2:0]}), .CI(1'b0), .SUM({N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, 
        N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47}) );
  ALU_N32_DW01_cmp6_5 r59 ( .A({DATA1[31:26], n60, DATA1[24:23], n49, 
        DATA1[21], n23, n29, DATA1[18:15], n56, n100, DATA1[12:11], n112, n110, 
        n114, n43, n5, n64, n52, n72, DATA1[2], n102, n107}), .B({DATA2[31:29], 
        n103, DATA2[27:18], n46, n116, n82, DATA2[14], n58, DATA2[12:10], n57, 
        n66, n53, DATA2[6:5], n81, n79, n119, DATA2[1], n101}), .TC(1'b1), 
        .LE(N111), .GE(N112) );
endmodule


module DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 ( CLK, RST, IR_IN, 
        IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
        RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
        EQ_COND, IS_JUMP, .ALU_OPCODE({\ALU_OPCODE[3] , \ALU_OPCODE[2] , 
        \ALU_OPCODE[1] , \ALU_OPCODE[0] }), JUMP_EN, PC_LATCH_EN, IS_JAL, 
        WB_MUX_SEL, RF_WE, D_ADDR, D_DATA_IN, D_DATA_OUT, PC_IN, PC_BUS );
  input [31:0] IR_IN;
  output [5:0] D_ADDR;
  output [31:0] D_DATA_IN;
  input [31:0] D_DATA_OUT;
  input [31:0] PC_IN;
  output [31:0] PC_BUS;
  input CLK, RST, IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN,
         RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN,
         EQ_COND, IS_JUMP, \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] ,
         \ALU_OPCODE[0] , JUMP_EN, PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE;
  wire   branch_taken, PC_MUX_SEL, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [3:0] ALU_OPCODE;
  wire   [31:0] current_PC1;
  wire   [31:0] current_PC2;
  wire   [31:0] current_PC3;
  wire   [31:0] current_PC4;
  wire   [31:0] next_NPC;
  wire   [31:0] current_NPC;
  wire   [25:0] current_IW;
  wire   [25:0] IMM_IN;
  wire   [4:0] WB1_IN;
  wire   [4:0] WB2_IN;
  wire   [4:0] WB2_OUT;
  wire   [4:0] WB3_OUT;
  wire   [31:0] next_ALU_OUT;
  wire   [31:6] current_ALU_OUT;
  wire   [31:0] B_OUT;
  wire   [31:0] current_ALU_OUT2;
  wire   [31:0] A_OUT;
  wire   [31:0] ALU_OP1;
  wire   [31:0] IMM_OUT;
  wire   [31:0] ALU_OP2;
  wire   [31:0] OUT_MUX_DATA;
  wire   [31:0] WB_DATA;
  wire   [4:0] WB_ADDR;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5;

  BUF_X1 U3 ( .A(D_ADDR[2]), .Z(n1) );
  BUF_X1 U4 ( .A(D_ADDR[0]), .Z(n2) );
  BUF_X1 U5 ( .A(D_ADDR[1]), .Z(n3) );
  BUF_X1 U6 ( .A(D_ADDR[3]), .Z(n4) );
  BUF_X1 U7 ( .A(D_ADDR[4]), .Z(n5) );
  BUF_X1 U8 ( .A(D_ADDR[5]), .Z(n6) );
  CLKBUF_X1 U9 ( .A(IS_JUMP), .Z(n7) );
  CLKBUF_X3 U10 ( .A(RST), .Z(n8) );
  REG_GENERIC_NBIT32_9 PC_REG ( .CLK(CLK), .RST(n8), .EN(PC_LATCH_EN), 
        .DATA_IN(PC_IN), .DATA_OUT(current_PC1) );
  REG_GENERIC_NBIT32_8 PC2_REG ( .CLK(CLK), .RST(n8), .EN(PC_LATCH_EN), 
        .DATA_IN(current_PC1), .DATA_OUT(current_PC2) );
  REG_GENERIC_NBIT32_7 PC3_REG ( .CLK(CLK), .RST(n8), .EN(PC_LATCH_EN), 
        .DATA_IN(current_PC2), .DATA_OUT(current_PC3) );
  REG_GENERIC_NBIT32_6 PC4_REG ( .CLK(CLK), .RST(n8), .EN(PC_LATCH_EN), 
        .DATA_IN(current_PC3), .DATA_OUT(current_PC4) );
  REG_GENERIC_NBIT32_5 NPC_REG ( .CLK(CLK), .RST(n8), .EN(NPC_LATCH_EN), 
        .DATA_IN(next_NPC), .DATA_OUT(current_NPC) );
  REG_GENERIC_NBIT32_4 IR_REG ( .CLK(CLK), .RST(n8), .EN(IR_LATCH_EN), 
        .DATA_IN(IR_IN), .DATA_OUT({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, current_IW}) );
  REG_GENERIC_NBIT26 IMM_REG ( .CLK(CLK), .RST(n8), .EN(RegIMM_LATCH_EN), 
        .DATA_IN(current_IW), .DATA_OUT(IMM_IN) );
  REG_GENERIC_NBIT5_0 WB1_REG ( .CLK(CLK), .RST(n8), .EN(1'b1), .DATA_IN(
        WB1_IN), .DATA_OUT(WB2_IN) );
  REG_GENERIC_NBIT5_2 WB2_REG ( .CLK(CLK), .RST(n8), .EN(ALU_OUTREG_EN), 
        .DATA_IN(WB2_IN), .DATA_OUT(WB2_OUT) );
  REG_GENERIC_NBIT5_1 WB3_REG ( .CLK(CLK), .RST(n8), .EN(1'b1), .DATA_IN(
        WB2_OUT), .DATA_OUT(WB3_OUT) );
  REG_GENERIC_NBIT32_3 ALU_OUT_REG ( .CLK(CLK), .RST(n8), .EN(ALU_OUTREG_EN), 
        .DATA_IN(next_ALU_OUT), .DATA_OUT({current_ALU_OUT, D_ADDR}) );
  REG_GENERIC_NBIT32_2 B_OUT_REG ( .CLK(CLK), .RST(n8), .EN(ALU_OUTREG_EN), 
        .DATA_IN(B_OUT), .DATA_OUT(D_DATA_IN) );
  REG_GENERIC_NBIT32_1 ALU_OUT_REG2 ( .CLK(CLK), .RST(n8), .EN(1'b1), 
        .DATA_IN({current_ALU_OUT, n6, n5, n4, n1, n3, n2}), .DATA_OUT(
        current_ALU_OUT2) );
  BRANCHING_UNIT_N32 BU ( .CLK(CLK), .RST(n8), .Reg_A(A_OUT), .EQ_cond(EQ_COND), .IS_JUMP(n7), .branch_taken(branch_taken) );
  MUX21_GENERIC_NBIT32_0 PC_MUX ( .A(current_NPC), .B({current_ALU_OUT, n6, n5, 
        n4, n1, n3, n2}), .SEL(PC_MUX_SEL), .Y(PC_BUS) );
  MUX21 J_MUX ( .A(1'b0), .B(branch_taken), .SEL(JUMP_EN), .Y(PC_MUX_SEL) );
  MUX21_GENERIC_NBIT5_0 RD_MUX ( .A(current_IW[15:11]), .B(current_IW[20:16]), 
        .SEL(RegIMM_LATCH_EN), .Y(WB1_IN) );
  MUX21_GENERIC_NBIT32_4 OP1_MUX ( .A(A_OUT), .B(current_PC2), .SEL(MUXA_SEL), 
        .Y(ALU_OP1) );
  MUX21_GENERIC_NBIT32_3 OP2_MUX ( .A(B_OUT), .B(IMM_OUT), .SEL(MUXB_SEL), .Y(
        ALU_OP2) );
  MUX21_GENERIC_NBIT32_2 OUT_MUX ( .A(D_DATA_OUT), .B(current_ALU_OUT2), .SEL(
        WB_MUX_SEL), .Y(OUT_MUX_DATA) );
  MUX21_GENERIC_NBIT32_1 JAL_DATA_MUX ( .A(OUT_MUX_DATA), .B(current_PC4), 
        .SEL(IS_JAL), .Y(WB_DATA) );
  MUX21_GENERIC_NBIT5_1 JAL_ADDR_MUX ( .A(WB3_OUT), .B({1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1}), .SEL(IS_JAL), .Y(WB_ADDR) );
  ADDER_N32 PC_ADDER ( .CURR_ADDR(PC_BUS), .NEXT_ADDR(next_NPC) );
  REGISTER_FILE_NBIT32_NREG32 RF ( .CLK(CLK), .RST(n8), .EN(1'b1), .RD1(
        RegA_LATCH_EN), .RD2(RegB_LATCH_EN), .WR(RF_WE), .ADD_WR(WB_ADDR), 
        .ADD_RD1(current_IW[25:21]), .ADD_RD2(current_IW[20:16]), .DATAIN(
        WB_DATA), .OUT1(A_OUT), .OUT2(B_OUT) );
  EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26 EXT ( .NOT_EXT_IMM(IMM_IN), .SIGNED_IMM(
        SIGNED_IMM), .IS_JUMP(IS_JUMP), .EXT_IMM(IMM_OUT) );
  ALU_N32 ALU_i ( .FUNC({\ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), .DATA1(ALU_OP1), .DATA2(ALU_OP2), .OUTALU(
        next_ALU_OUT) );
endmodule


module dlx_cu ( Clk, Rst, IR_IN, IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, 
        RegB_LATCH_EN, RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, 
        ALU_OUTREG_EN, EQ_COND, IS_JUMP, .ALU_OPCODE({\ALU_OPCODE[3] , 
        \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] }), DRAM_WE, 
        LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE );
  input [31:0] IR_IN;
  input Clk, Rst;
  output IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN,
         RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN,
         EQ_COND, IS_JUMP, \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] ,
         \ALU_OPCODE[0] , DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, IS_JAL,
         WB_MUX_SEL, RF_WE;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26, n34, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83;
  wire   [3:0] ALU_OPCODE;
  wire   [17:0] cw;
  wire   [15:0] cw1;
  wire   [12:0] cw2;
  wire   [6:0] cw3;
  wire   [2:0] cw4;
  wire   [3:0] aluOpcode1;
  wire   [3:0] aluOpcode2;
  wire   [3:0] aluOpcode_i;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];

  DFFS_X1 \cw1_reg[17]  ( .D(cw[17]), .CK(Clk), .SN(Rst), .Q(IR_LATCH_EN) );
  DFFS_X1 \cw1_reg[16]  ( .D(cw[17]), .CK(Clk), .SN(Rst), .Q(NPC_LATCH_EN) );
  DFFR_X1 \cw1_reg[15]  ( .D(cw[9]), .CK(Clk), .RN(Rst), .Q(cw1[15]) );
  DFFR_X1 \cw2_reg[15]  ( .D(cw1[15]), .CK(Clk), .RN(Rst), .Q(RegA_LATCH_EN)
         );
  DFFR_X1 \cw1_reg[14]  ( .D(cw[14]), .CK(Clk), .RN(Rst), .Q(cw1[14]) );
  DFFR_X1 \cw2_reg[14]  ( .D(cw1[14]), .CK(Clk), .RN(Rst), .Q(RegB_LATCH_EN)
         );
  DFFR_X1 \cw1_reg[13]  ( .D(cw[13]), .CK(Clk), .RN(Rst), .Q(cw1[13]) );
  DFFR_X1 \cw2_reg[13]  ( .D(cw1[13]), .CK(Clk), .RN(Rst), .Q(RegIMM_LATCH_EN)
         );
  DFFR_X1 \cw1_reg[12]  ( .D(cw[12]), .CK(Clk), .RN(Rst), .Q(cw1[12]) );
  DFFR_X1 \cw2_reg[12]  ( .D(cw1[12]), .CK(Clk), .RN(Rst), .Q(cw2[12]) );
  DFFR_X1 \cw1_reg[11]  ( .D(cw[4]), .CK(Clk), .RN(Rst), .Q(cw1[11]) );
  DFFR_X1 \cw2_reg[11]  ( .D(cw1[11]), .CK(Clk), .RN(Rst), .Q(cw2[11]) );
  DFFR_X1 \cw1_reg[10]  ( .D(cw[13]), .CK(Clk), .RN(Rst), .Q(cw1[10]) );
  DFFR_X1 \cw2_reg[10]  ( .D(cw1[10]), .CK(Clk), .RN(Rst), .Q(cw2[10]) );
  DFFR_X1 \cw1_reg[9]  ( .D(cw[9]), .CK(Clk), .RN(Rst), .Q(cw1[9]) );
  DFFR_X1 \cw2_reg[9]  ( .D(cw1[9]), .CK(Clk), .RN(Rst), .Q(cw2[9]) );
  DFFR_X1 \cw1_reg[8]  ( .D(cw[8]), .CK(Clk), .RN(Rst), .Q(cw1[8]) );
  DFFR_X1 \cw2_reg[8]  ( .D(cw1[8]), .CK(Clk), .RN(Rst), .Q(cw2[8]) );
  DFFR_X1 \cw1_reg[7]  ( .D(n83), .CK(Clk), .RN(Rst), .Q(cw1[7]) );
  DFFR_X1 \cw2_reg[7]  ( .D(cw1[7]), .CK(Clk), .RN(Rst), .Q(cw2[7]) );
  DFFR_X1 \cw1_reg[6]  ( .D(cw[6]), .CK(Clk), .RN(Rst), .Q(cw1[6]) );
  DFFR_X1 \cw2_reg[6]  ( .D(cw1[6]), .CK(Clk), .RN(Rst), .Q(cw2[6]) );
  DFFR_X1 \cw1_reg[5]  ( .D(cw[5]), .CK(Clk), .RN(Rst), .Q(cw1[5]) );
  DFFR_X1 \cw2_reg[5]  ( .D(cw1[5]), .CK(Clk), .RN(Rst), .Q(cw2[5]) );
  DFFR_X1 \cw1_reg[4]  ( .D(cw[4]), .CK(Clk), .RN(Rst), .Q(cw1[4]) );
  DFFR_X1 \cw2_reg[4]  ( .D(cw1[4]), .CK(Clk), .RN(Rst), .Q(cw2[4]) );
  DFFS_X1 \cw1_reg[3]  ( .D(cw[3]), .CK(Clk), .SN(Rst), .Q(cw1[3]) );
  DFFS_X1 \cw2_reg[3]  ( .D(cw1[3]), .CK(Clk), .SN(Rst), .Q(cw2[3]) );
  SDFFR_X1 \cw1_reg[2]  ( .D(1'b0), .SI(n83), .SE(IR_IN_26), .CK(Clk), .RN(Rst), .Q(cw1[2]) );
  DFFR_X1 \cw2_reg[2]  ( .D(cw1[2]), .CK(Clk), .RN(Rst), .Q(cw2[2]) );
  DFFR_X1 \cw1_reg[1]  ( .D(cw[1]), .CK(Clk), .RN(Rst), .Q(cw1[1]) );
  DFFR_X1 \cw2_reg[1]  ( .D(cw1[1]), .CK(Clk), .RN(Rst), .Q(cw2[1]) );
  SDFFR_X1 \cw1_reg[0]  ( .D(1'b1), .SI(cw[1]), .SE(n34), .CK(Clk), .RN(Rst), 
        .Q(cw1[0]) );
  DFFR_X1 \cw2_reg[0]  ( .D(cw1[0]), .CK(Clk), .RN(Rst), .Q(cw2[0]) );
  DFFR_X1 \cw3_reg[12]  ( .D(cw2[12]), .CK(Clk), .RN(Rst), .Q(SIGNED_IMM) );
  DFFR_X1 \cw3_reg[11]  ( .D(cw2[11]), .CK(Clk), .RN(Rst), .Q(MUXA_SEL) );
  DFFR_X1 \cw3_reg[10]  ( .D(cw2[10]), .CK(Clk), .RN(Rst), .Q(MUXB_SEL) );
  DFFR_X1 \cw3_reg[9]  ( .D(cw2[9]), .CK(Clk), .RN(Rst), .Q(ALU_OUTREG_EN) );
  DFFR_X1 \cw3_reg[8]  ( .D(cw2[8]), .CK(Clk), .RN(Rst), .Q(EQ_COND) );
  DFFR_X1 \cw3_reg[6]  ( .D(cw2[6]), .CK(Clk), .RN(Rst), .Q(cw3[6]) );
  DFFR_X1 \cw3_reg[5]  ( .D(cw2[5]), .CK(Clk), .RN(Rst), .Q(cw3[5]) );
  DFFR_X1 \cw3_reg[4]  ( .D(cw2[4]), .CK(Clk), .RN(Rst), .Q(cw3[4]) );
  DFFS_X1 \cw3_reg[3]  ( .D(cw2[3]), .CK(Clk), .SN(Rst), .Q(cw3[3]) );
  DFFR_X1 \cw3_reg[2]  ( .D(cw2[2]), .CK(Clk), .RN(Rst), .Q(cw3[2]) );
  DFFR_X1 \cw3_reg[1]  ( .D(cw2[1]), .CK(Clk), .RN(Rst), .Q(cw3[1]) );
  DFFR_X1 \cw3_reg[0]  ( .D(cw2[0]), .CK(Clk), .RN(Rst), .Q(cw3[0]) );
  DFFR_X1 \cw4_reg[6]  ( .D(cw3[6]), .CK(Clk), .RN(Rst), .Q(DRAM_WE) );
  DFFR_X1 \cw4_reg[5]  ( .D(cw3[5]), .CK(Clk), .RN(Rst), .Q(LMD_LATCH_EN) );
  DFFR_X1 \cw4_reg[4]  ( .D(cw3[4]), .CK(Clk), .RN(Rst), .Q(JUMP_EN) );
  DFFS_X1 \cw4_reg[3]  ( .D(cw3[3]), .CK(Clk), .SN(Rst), .Q(PC_LATCH_EN) );
  DFFR_X1 \cw4_reg[2]  ( .D(cw3[2]), .CK(Clk), .RN(Rst), .Q(cw4[2]) );
  DFFR_X1 \cw4_reg[1]  ( .D(cw3[1]), .CK(Clk), .RN(Rst), .Q(cw4[1]) );
  DFFR_X1 \cw4_reg[0]  ( .D(cw3[0]), .CK(Clk), .RN(Rst), .Q(cw4[0]) );
  DFFR_X1 \cw5_reg[2]  ( .D(cw4[2]), .CK(Clk), .RN(Rst), .Q(IS_JAL) );
  DFFR_X1 \cw5_reg[1]  ( .D(cw4[1]), .CK(Clk), .RN(Rst), .Q(WB_MUX_SEL) );
  DFFR_X1 \cw5_reg[0]  ( .D(cw4[0]), .CK(Clk), .RN(Rst), .Q(RF_WE) );
  DFFR_X1 \aluOpcode1_reg[3]  ( .D(aluOpcode_i[3]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[3]) );
  DFFR_X1 \aluOpcode1_reg[2]  ( .D(aluOpcode_i[2]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[2]) );
  DFFR_X1 \aluOpcode1_reg[1]  ( .D(aluOpcode_i[1]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[1]) );
  DFFR_X1 \aluOpcode1_reg[0]  ( .D(aluOpcode_i[0]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[0]) );
  DFFR_X1 \aluOpcode2_reg[3]  ( .D(aluOpcode1[3]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[3]) );
  DFFR_X1 \aluOpcode3_reg[3]  ( .D(aluOpcode2[3]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[3]) );
  DFFR_X1 \aluOpcode2_reg[2]  ( .D(aluOpcode1[2]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[2]) );
  DFFR_X1 \aluOpcode3_reg[2]  ( .D(aluOpcode2[2]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[2]) );
  DFFR_X1 \aluOpcode2_reg[1]  ( .D(aluOpcode1[1]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[1]) );
  DFFR_X1 \aluOpcode3_reg[1]  ( .D(aluOpcode2[1]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[1]) );
  DFFR_X1 \aluOpcode2_reg[0]  ( .D(aluOpcode1[0]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[0]) );
  DFFR_X1 \aluOpcode3_reg[0]  ( .D(aluOpcode2[0]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[0]) );
  DFFR_X1 \cw3_reg[7]  ( .D(cw2[7]), .CK(Clk), .RN(Rst), .Q(IS_JUMP) );
  INV_X1 U5 ( .A(n42), .ZN(n29) );
  NOR2_X1 U6 ( .A1(n78), .A2(n59), .ZN(n26) );
  AND2_X1 U7 ( .A1(n22), .A2(n53), .ZN(n3) );
  AND2_X1 U8 ( .A1(n65), .A2(n76), .ZN(n4) );
  AND2_X1 U9 ( .A1(n7), .A2(n68), .ZN(n5) );
  NAND4_X1 U10 ( .A1(n33), .A2(n32), .A3(n31), .A4(n30), .ZN(aluOpcode_i[0])
         );
  NOR2_X1 U11 ( .A1(cw[4]), .A2(n29), .ZN(n30) );
  NOR2_X1 U12 ( .A1(n17), .A2(n11), .ZN(n33) );
  AOI22_X1 U13 ( .A1(n28), .A2(n27), .B1(n26), .B2(n25), .ZN(n31) );
  AND3_X1 U14 ( .A1(n5), .A2(n34), .A3(n72), .ZN(n6) );
  AND3_X1 U15 ( .A1(n60), .A2(n59), .A3(n58), .ZN(n7) );
  OAI22_X1 U16 ( .A1(n8), .A2(n60), .B1(IR_IN_30), .B2(n68), .ZN(n17) );
  AND2_X1 U17 ( .A1(IR_IN_27), .A2(n77), .ZN(n8) );
  OAI21_X1 U18 ( .B1(IR_IN[1]), .B2(n51), .A(n43), .ZN(n27) );
  AND2_X1 U19 ( .A1(IR_IN_28), .A2(n78), .ZN(n9) );
  AND2_X1 U20 ( .A1(IR_IN_30), .A2(IR_IN_26), .ZN(n10) );
  NAND2_X1 U21 ( .A1(n23), .A2(IR_IN[0]), .ZN(n32) );
  INV_X1 U22 ( .A(n47), .ZN(n23) );
  AND2_X1 U23 ( .A1(IR_IN[1]), .A2(n37), .ZN(n11) );
  INV_X1 U24 ( .A(IR_IN_27), .ZN(n78) );
  INV_X1 U25 ( .A(IR_IN_31), .ZN(n25) );
  NAND2_X1 U26 ( .A1(n9), .A2(n25), .ZN(n82) );
  INV_X1 U27 ( .A(n82), .ZN(n66) );
  INV_X1 U28 ( .A(IR_IN_30), .ZN(n65) );
  INV_X1 U29 ( .A(IR_IN_29), .ZN(n24) );
  NAND2_X1 U30 ( .A1(n65), .A2(n24), .ZN(n35) );
  INV_X1 U31 ( .A(n35), .ZN(n79) );
  NAND2_X1 U32 ( .A1(n66), .A2(n79), .ZN(n63) );
  INV_X1 U33 ( .A(IR_IN_28), .ZN(n77) );
  NAND3_X1 U34 ( .A1(n79), .A2(n8), .A3(n25), .ZN(n80) );
  NAND2_X1 U35 ( .A1(n63), .A2(n80), .ZN(cw[4]) );
  INV_X1 U36 ( .A(IR_IN_26), .ZN(n76) );
  NAND3_X1 U37 ( .A1(n4), .A2(IR_IN_29), .A3(n25), .ZN(n60) );
  NAND3_X1 U38 ( .A1(IR_IN_26), .A2(IR_IN_31), .A3(n8), .ZN(n68) );
  INV_X1 U39 ( .A(IR_IN[0]), .ZN(n50) );
  INV_X1 U40 ( .A(IR_IN[3]), .ZN(n49) );
  NAND2_X1 U41 ( .A1(n50), .A2(n49), .ZN(n44) );
  INV_X1 U42 ( .A(n44), .ZN(n28) );
  INV_X1 U43 ( .A(IR_IN[5]), .ZN(n16) );
  OR3_X1 U44 ( .A1(IR_IN[6]), .A2(IR_IN[7]), .A3(IR_IN[4]), .ZN(n12) );
  OR4_X1 U45 ( .A1(IR_IN[9]), .A2(IR_IN[10]), .A3(IR_IN[8]), .A4(n12), .ZN(n18) );
  NAND3_X1 U46 ( .A1(n4), .A2(n25), .A3(n77), .ZN(n72) );
  INV_X1 U47 ( .A(n72), .ZN(n13) );
  NAND2_X1 U48 ( .A1(n13), .A2(n78), .ZN(n61) );
  INV_X1 U49 ( .A(n61), .ZN(n14) );
  NAND2_X1 U50 ( .A1(n14), .A2(n24), .ZN(n75) );
  INV_X1 U51 ( .A(IR_IN[2]), .ZN(n54) );
  NOR3_X1 U52 ( .A1(n18), .A2(n75), .A3(n54), .ZN(n15) );
  NAND3_X1 U53 ( .A1(n28), .A2(n16), .A3(n15), .ZN(n55) );
  INV_X1 U54 ( .A(n55), .ZN(n37) );
  INV_X1 U55 ( .A(n75), .ZN(n20) );
  INV_X1 U56 ( .A(n18), .ZN(n19) );
  NAND3_X1 U57 ( .A1(IR_IN[5]), .A2(n20), .A3(n19), .ZN(n51) );
  INV_X1 U58 ( .A(n51), .ZN(n21) );
  NAND2_X1 U59 ( .A1(n21), .A2(IR_IN[2]), .ZN(n43) );
  INV_X1 U60 ( .A(n43), .ZN(n22) );
  INV_X1 U61 ( .A(IR_IN[1]), .ZN(n53) );
  NAND2_X1 U62 ( .A1(n3), .A2(IR_IN[3]), .ZN(n47) );
  NAND4_X1 U63 ( .A1(IR_IN_30), .A2(IR_IN_28), .A3(n24), .A4(n76), .ZN(n59) );
  NAND2_X1 U64 ( .A1(n66), .A2(IR_IN_29), .ZN(n62) );
  INV_X1 U65 ( .A(n62), .ZN(n64) );
  NAND2_X1 U66 ( .A1(n64), .A2(n10), .ZN(n42) );
  NAND3_X1 U67 ( .A1(n66), .A2(n35), .A3(n76), .ZN(n41) );
  INV_X1 U68 ( .A(n60), .ZN(n39) );
  NOR3_X1 U69 ( .A1(IR_IN[2]), .A2(n44), .A3(n51), .ZN(n36) );
  MUX2_X1 U70 ( .A(n37), .B(n36), .S(IR_IN[1]), .Z(n38) );
  AOI221_X1 U71 ( .B1(n3), .B2(n50), .C1(n39), .C2(n8), .A(n38), .ZN(n40) );
  NAND4_X1 U72 ( .A1(n42), .A2(n47), .A3(n41), .A4(n40), .ZN(aluOpcode_i[1])
         );
  OAI33_X1 U73 ( .A1(n60), .A2(n77), .A3(n78), .B1(n44), .B2(n43), .B3(n53), 
        .ZN(n45) );
  AOI21_X1 U74 ( .B1(n3), .B2(IR_IN[0]), .A(n45), .ZN(n46) );
  OAI211_X1 U75 ( .C1(n4), .C2(n62), .A(n47), .B(n46), .ZN(aluOpcode_i[2]) );
  NAND3_X1 U76 ( .A1(IR_IN_29), .A2(n10), .A3(n78), .ZN(n58) );
  INV_X1 U77 ( .A(n58), .ZN(n69) );
  INV_X1 U78 ( .A(n59), .ZN(n48) );
  AOI21_X1 U79 ( .B1(n69), .B2(n77), .A(n48), .ZN(n57) );
  NOR3_X1 U80 ( .A1(n51), .A2(n50), .A3(n49), .ZN(n52) );
  NAND3_X1 U81 ( .A1(n54), .A2(n53), .A3(n52), .ZN(n56) );
  OAI211_X1 U82 ( .C1(IR_IN_31), .C2(n57), .A(n56), .B(n55), .ZN(
        aluOpcode_i[3]) );
  NAND3_X1 U83 ( .A1(n7), .A2(n62), .A3(n61), .ZN(cw[1]) );
  NAND3_X1 U84 ( .A1(n79), .A2(IR_IN_26), .A3(n8), .ZN(n34) );
  INV_X1 U85 ( .A(n80), .ZN(n83) );
  NAND2_X1 U86 ( .A1(n82), .A2(n6), .ZN(cw[3]) );
  NOR2_X1 U87 ( .A1(IR_IN_29), .A2(n68), .ZN(cw[5]) );
  NAND4_X1 U88 ( .A1(IR_IN_29), .A2(IR_IN_31), .A3(IR_IN_27), .A4(IR_IN_26), 
        .ZN(n74) );
  INV_X1 U89 ( .A(n74), .ZN(cw[6]) );
  OAI21_X1 U90 ( .B1(IR_IN_26), .B2(n63), .A(n80), .ZN(cw[8]) );
  OAI21_X1 U91 ( .B1(n10), .B2(n82), .A(n6), .ZN(cw[9]) );
  AOI21_X1 U92 ( .B1(n66), .B2(n65), .A(n64), .ZN(n67) );
  NAND3_X1 U93 ( .A1(n5), .A2(n80), .A3(n67), .ZN(cw[13]) );
  NAND3_X1 U94 ( .A1(IR_IN_29), .A2(IR_IN_30), .A3(n9), .ZN(n73) );
  INV_X1 U95 ( .A(n68), .ZN(n70) );
  NOR3_X1 U96 ( .A1(n70), .A2(cw[4]), .A3(n69), .ZN(n71) );
  NAND3_X1 U97 ( .A1(n73), .A2(n72), .A3(n71), .ZN(cw[12]) );
  NAND2_X1 U98 ( .A1(n75), .A2(n74), .ZN(cw[14]) );
  NAND4_X1 U99 ( .A1(n79), .A2(n78), .A3(n77), .A4(n76), .ZN(n81) );
  NAND4_X1 U100 ( .A1(n5), .A2(n82), .A3(n81), .A4(n80), .ZN(cw[17]) );
endmodule


module DLX ( CLK, RST, I_ADDR, I_DATA, D_RR, D_WR, D_ADDR, D_DATA_IN, 
        D_DATA_OUT );
  output [31:0] I_ADDR;
  input [31:0] I_DATA;
  output [5:0] D_ADDR;
  output [31:0] D_DATA_IN;
  input [31:0] D_DATA_OUT;
  input CLK, RST;
  output D_RR, D_WR;
  wire   PC_LATCH_EN, IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN,
         RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN,
         EQ_COND, IS_JUMP, JUMP_EN, IS_JAL, WB_MUX_SEL, RF_WE, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [31:0] PC_BUS;
  wire   [3:0] ALU_OPCODE;

  BUF_X1 U1 ( .A(I_ADDR[3]), .Z(n1) );
  BUF_X1 U2 ( .A(I_ADDR[22]), .Z(n2) );
  BUF_X1 U3 ( .A(I_ADDR[25]), .Z(n3) );
  BUF_X1 U4 ( .A(I_ADDR[4]), .Z(n4) );
  BUF_X1 U5 ( .A(I_ADDR[6]), .Z(n5) );
  BUF_X1 U6 ( .A(I_ADDR[7]), .Z(n6) );
  BUF_X1 U7 ( .A(I_ADDR[9]), .Z(n7) );
  BUF_X1 U8 ( .A(I_ADDR[10]), .Z(n8) );
  BUF_X1 U9 ( .A(I_ADDR[14]), .Z(n9) );
  BUF_X1 U10 ( .A(I_ADDR[15]), .Z(n10) );
  BUF_X1 U11 ( .A(I_ADDR[18]), .Z(n11) );
  BUF_X1 U12 ( .A(I_ADDR[20]), .Z(n12) );
  BUF_X1 U13 ( .A(I_ADDR[23]), .Z(n13) );
  BUF_X1 U14 ( .A(I_ADDR[26]), .Z(n14) );
  BUF_X1 U15 ( .A(I_ADDR[27]), .Z(n15) );
  BUF_X1 U16 ( .A(I_ADDR[28]), .Z(n16) );
  BUF_X1 U17 ( .A(I_ADDR[30]), .Z(n17) );
  CLKBUF_X1 U18 ( .A(I_ADDR[0]), .Z(n18) );
  CLKBUF_X1 U19 ( .A(I_ADDR[1]), .Z(n19) );
  CLKBUF_X1 U20 ( .A(I_ADDR[2]), .Z(n20) );
  CLKBUF_X1 U21 ( .A(I_ADDR[8]), .Z(n21) );
  CLKBUF_X1 U22 ( .A(I_ADDR[11]), .Z(n22) );
  CLKBUF_X1 U23 ( .A(I_ADDR[12]), .Z(n23) );
  CLKBUF_X1 U24 ( .A(I_ADDR[13]), .Z(n24) );
  CLKBUF_X1 U25 ( .A(I_ADDR[17]), .Z(n25) );
  CLKBUF_X1 U26 ( .A(I_ADDR[19]), .Z(n26) );
  CLKBUF_X1 U27 ( .A(I_ADDR[31]), .Z(n27) );
  REG_GENERIC_NBIT32_0 PC_REG ( .CLK(CLK), .RST(RST), .EN(PC_LATCH_EN), 
        .DATA_IN(PC_BUS), .DATA_OUT(I_ADDR) );
  DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 DP ( .CLK(CLK), .RST(RST), 
        .IR_IN(I_DATA), .IR_LATCH_EN(IR_LATCH_EN), .NPC_LATCH_EN(NPC_LATCH_EN), 
        .RegA_LATCH_EN(RegA_LATCH_EN), .RegB_LATCH_EN(RegB_LATCH_EN), 
        .RegIMM_LATCH_EN(RegIMM_LATCH_EN), .SIGNED_IMM(SIGNED_IMM), .MUXA_SEL(
        MUXA_SEL), .MUXB_SEL(MUXB_SEL), .ALU_OUTREG_EN(ALU_OUTREG_EN), 
        .EQ_COND(EQ_COND), .IS_JUMP(IS_JUMP), .ALU_OPCODE(ALU_OPCODE), 
        .JUMP_EN(JUMP_EN), .PC_LATCH_EN(PC_LATCH_EN), .IS_JAL(IS_JAL), 
        .WB_MUX_SEL(WB_MUX_SEL), .RF_WE(RF_WE), .D_ADDR(D_ADDR), .D_DATA_IN(
        D_DATA_IN), .D_DATA_OUT(D_DATA_OUT), .PC_IN({n27, n17, I_ADDR[29], n16, 
        n15, n14, n3, I_ADDR[24], n13, n2, I_ADDR[21], n12, n26, n11, n25, 
        I_ADDR[16], n10, n9, n24, n23, n22, n8, n7, n21, n6, n5, I_ADDR[5], n4, 
        n1, n20, n19, n18}), .PC_BUS(PC_BUS) );
  dlx_cu CU ( .Clk(CLK), .Rst(RST), .IR_IN(I_DATA), .IR_LATCH_EN(IR_LATCH_EN), 
        .NPC_LATCH_EN(NPC_LATCH_EN), .RegA_LATCH_EN(RegA_LATCH_EN), 
        .RegB_LATCH_EN(RegB_LATCH_EN), .RegIMM_LATCH_EN(RegIMM_LATCH_EN), 
        .SIGNED_IMM(SIGNED_IMM), .MUXA_SEL(MUXA_SEL), .MUXB_SEL(MUXB_SEL), 
        .ALU_OUTREG_EN(ALU_OUTREG_EN), .EQ_COND(EQ_COND), .IS_JUMP(IS_JUMP), 
        .ALU_OPCODE(ALU_OPCODE), .DRAM_WE(D_WR), .LMD_LATCH_EN(D_RR), 
        .JUMP_EN(JUMP_EN), .PC_LATCH_EN(PC_LATCH_EN), .IS_JAL(IS_JAL), 
        .WB_MUX_SEL(WB_MUX_SEL), .RF_WE(RF_WE) );
endmodule

