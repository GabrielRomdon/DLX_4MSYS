
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOpType is (NOP, ADDS, SUBS, ANDS, ORS, XORS, SLE, SGE, SNE, SRLS, SLLS)
   ;
attribute ENUM_ENCODING of aluOpType : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOpType(arg : in std_logic_vector( 1 to 4 )) 
               return aluOpType;
   function aluOpType_to_std_logic_vector(arg : in aluOpType) return 
               std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOpType(arg : in std_logic_vector( 1 to 4 )) 
   return aluOpType is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "0000" => return NOP;
         when "0001" => return ADDS;
         when "0010" => return SUBS;
         when "0011" => return ANDS;
         when "0100" => return ORS;
         when "0101" => return XORS;
         when "0110" => return SLE;
         when "0111" => return SGE;
         when "1000" => return SNE;
         when "1001" => return SRLS;
         when "1010" => return SLLS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOpType_to_std_logic_vector(arg : in aluOpType) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "0000";
         when ADDS => return "0001";
         when SUBS => return "0010";
         when ANDS => return "0011";
         when ORS => return "0100";
         when XORS => return "0101";
         when SLE => return "0110";
         when SGE => return "0111";
         when SNE => return "1000";
         when SRLS => return "1001";
         when SLLS => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_N32_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end ADDER_N32_DW01_add_0;

architecture SYN_rpl of ADDER_N32_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, SUM_3_port,
      SUM_4_port, SUM_5_port, SUM_6_port, SUM_7_port, SUM_8_port, SUM_9_port, 
      SUM_10_port, SUM_11_port, SUM_12_port, SUM_13_port, SUM_14_port, 
      SUM_15_port, SUM_16_port, SUM_17_port, SUM_18_port, SUM_19_port, 
      SUM_20_port, SUM_21_port, SUM_22_port, SUM_23_port, SUM_24_port, 
      SUM_25_port, SUM_26_port, SUM_27_port, SUM_28_port, SUM_29_port, 
      SUM_30_port, SUM_31_port, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n1);
   U2 : AND2_X1 port map( A1 => A(4), A2 => n1, ZN => n2);
   U3 : AND2_X1 port map( A1 => A(5), A2 => n2, ZN => n3);
   U4 : AND2_X1 port map( A1 => A(6), A2 => n3, ZN => n4);
   U5 : AND2_X1 port map( A1 => A(7), A2 => n4, ZN => n5);
   U6 : AND2_X1 port map( A1 => A(8), A2 => n5, ZN => n6);
   U7 : AND2_X1 port map( A1 => A(9), A2 => n6, ZN => n7);
   U8 : AND2_X1 port map( A1 => A(10), A2 => n7, ZN => n8);
   U9 : AND2_X1 port map( A1 => A(11), A2 => n8, ZN => n9);
   U10 : AND2_X1 port map( A1 => A(12), A2 => n9, ZN => n10);
   U11 : AND2_X1 port map( A1 => A(13), A2 => n10, ZN => n11);
   U12 : AND2_X1 port map( A1 => A(14), A2 => n11, ZN => n12);
   U13 : AND2_X1 port map( A1 => A(15), A2 => n12, ZN => n13);
   U14 : AND2_X1 port map( A1 => A(16), A2 => n13, ZN => n14);
   U15 : AND2_X1 port map( A1 => A(17), A2 => n14, ZN => n15);
   U16 : AND2_X1 port map( A1 => A(18), A2 => n15, ZN => n16);
   U17 : AND2_X1 port map( A1 => A(19), A2 => n16, ZN => n17);
   U18 : AND2_X1 port map( A1 => A(20), A2 => n17, ZN => n18);
   U19 : AND2_X1 port map( A1 => A(21), A2 => n18, ZN => n19);
   U20 : AND2_X1 port map( A1 => A(22), A2 => n19, ZN => n20);
   U21 : AND2_X1 port map( A1 => A(23), A2 => n20, ZN => n21);
   U22 : AND2_X1 port map( A1 => A(24), A2 => n21, ZN => n22);
   U23 : AND2_X1 port map( A1 => A(25), A2 => n22, ZN => n23);
   U24 : AND2_X1 port map( A1 => A(26), A2 => n23, ZN => n24);
   U25 : AND2_X1 port map( A1 => A(27), A2 => n24, ZN => n25);
   U26 : AND2_X1 port map( A1 => A(28), A2 => n25, ZN => n26);
   U27 : AND2_X1 port map( A1 => A(29), A2 => n26, ZN => n27);
   U28 : AND2_X1 port map( A1 => A(30), A2 => n27, ZN => n28);
   U29 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U30 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U31 : XOR2_X1 port map( A => A(4), B => n1, Z => SUM_4_port);
   U32 : XOR2_X1 port map( A => A(5), B => n2, Z => SUM_5_port);
   U33 : XOR2_X1 port map( A => A(6), B => n3, Z => SUM_6_port);
   U34 : XOR2_X1 port map( A => A(7), B => n4, Z => SUM_7_port);
   U35 : XOR2_X1 port map( A => A(8), B => n5, Z => SUM_8_port);
   U36 : XOR2_X1 port map( A => A(9), B => n6, Z => SUM_9_port);
   U37 : XOR2_X1 port map( A => A(10), B => n7, Z => SUM_10_port);
   U38 : XOR2_X1 port map( A => A(11), B => n8, Z => SUM_11_port);
   U39 : XOR2_X1 port map( A => A(12), B => n9, Z => SUM_12_port);
   U40 : XOR2_X1 port map( A => A(13), B => n10, Z => SUM_13_port);
   U41 : XOR2_X1 port map( A => A(14), B => n11, Z => SUM_14_port);
   U42 : XOR2_X1 port map( A => A(15), B => n12, Z => SUM_15_port);
   U43 : XOR2_X1 port map( A => A(16), B => n13, Z => SUM_16_port);
   U44 : XOR2_X1 port map( A => A(17), B => n14, Z => SUM_17_port);
   U45 : XOR2_X1 port map( A => A(18), B => n15, Z => SUM_18_port);
   U46 : XOR2_X1 port map( A => A(19), B => n16, Z => SUM_19_port);
   U47 : XOR2_X1 port map( A => A(20), B => n17, Z => SUM_20_port);
   U48 : XOR2_X1 port map( A => A(21), B => n18, Z => SUM_21_port);
   U49 : XOR2_X1 port map( A => A(22), B => n19, Z => SUM_22_port);
   U50 : XOR2_X1 port map( A => A(23), B => n20, Z => SUM_23_port);
   U51 : XOR2_X1 port map( A => A(24), B => n21, Z => SUM_24_port);
   U52 : XOR2_X1 port map( A => A(25), B => n22, Z => SUM_25_port);
   U53 : XOR2_X1 port map( A => A(26), B => n23, Z => SUM_26_port);
   U54 : XOR2_X1 port map( A => A(27), B => n24, Z => SUM_27_port);
   U55 : XOR2_X1 port map( A => A(28), B => n25, Z => SUM_28_port);
   U56 : XOR2_X1 port map( A => A(29), B => n26, Z => SUM_29_port);
   U57 : XOR2_X1 port map( A => A(30), B => n27, Z => SUM_30_port);
   U58 : XOR2_X1 port map( A => A(31), B => n28, Z => SUM_31_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end ALU_N32_DW01_cmp6_0;

architecture SYN_rpl of ALU_N32_DW01_cmp6_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal LE_port, GE_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208 : 
      std_logic;

begin
   LE <= LE_port;
   GE <= GE_port;
   
   U1 : INV_X1 port map( A => n135, ZN => n27);
   U2 : INV_X1 port map( A => n125, ZN => n23);
   U3 : INV_X1 port map( A => n115, ZN => n19);
   U4 : INV_X1 port map( A => n85, ZN => n7);
   U5 : INV_X1 port map( A => n105, ZN => n15);
   U6 : INV_X1 port map( A => n95, ZN => n11);
   U7 : INV_X1 port map( A => n131, ZN => n28);
   U8 : INV_X1 port map( A => n121, ZN => n24);
   U9 : INV_X1 port map( A => n111, ZN => n20);
   U10 : INV_X1 port map( A => n101, ZN => n16);
   U11 : INV_X1 port map( A => n91, ZN => n12);
   U12 : INV_X1 port map( A => n81, ZN => n8);
   U13 : INV_X1 port map( A => n140, ZN => n31);
   U14 : INV_X1 port map( A => n130, ZN => n26);
   U15 : INV_X1 port map( A => n114, ZN => n21);
   U16 : INV_X1 port map( A => n100, ZN => n14);
   U17 : INV_X1 port map( A => n84, ZN => n9);
   U18 : INV_X1 port map( A => n134, ZN => n29);
   U19 : INV_X1 port map( A => n104, ZN => n17);
   U20 : INV_X1 port map( A => n120, ZN => n22);
   U21 : INV_X1 port map( A => n90, ZN => n10);
   U22 : INV_X1 port map( A => n75, ZN => n5);
   U23 : INV_X1 port map( A => n139, ZN => n30);
   U24 : INV_X1 port map( A => n110, ZN => n18);
   U25 : INV_X1 port map( A => n80, ZN => n6);
   U26 : INV_X1 port map( A => n124, ZN => n25);
   U27 : INV_X1 port map( A => n94, ZN => n13);
   U28 : INV_X1 port map( A => B(2), ZN => n63);
   U29 : INV_X1 port map( A => B(0), ZN => n64);
   U30 : INV_X1 port map( A => n206, ZN => n32);
   U31 : INV_X1 port map( A => n65, ZN => LE_port);
   U32 : INV_X1 port map( A => A(31), ZN => n3);
   U33 : INV_X1 port map( A => A(1), ZN => n33);
   U34 : INV_X1 port map( A => n144, ZN => n34);
   U35 : INV_X1 port map( A => B(3), ZN => n62);
   U36 : INV_X1 port map( A => A(30), ZN => n4);
   U37 : INV_X1 port map( A => B(4), ZN => n61);
   U38 : INV_X1 port map( A => B(6), ZN => n59);
   U39 : INV_X1 port map( A => B(10), ZN => n55);
   U40 : INV_X1 port map( A => B(14), ZN => n51);
   U41 : INV_X1 port map( A => B(18), ZN => n47);
   U42 : INV_X1 port map( A => B(22), ZN => n43);
   U43 : INV_X1 port map( A => B(26), ZN => n39);
   U44 : INV_X1 port map( A => B(30), ZN => n35);
   U45 : INV_X1 port map( A => B(8), ZN => n57);
   U46 : INV_X1 port map( A => B(12), ZN => n53);
   U47 : INV_X1 port map( A => B(5), ZN => n60);
   U48 : INV_X1 port map( A => B(16), ZN => n49);
   U49 : INV_X1 port map( A => B(9), ZN => n56);
   U50 : INV_X1 port map( A => B(13), ZN => n52);
   U51 : INV_X1 port map( A => B(20), ZN => n45);
   U52 : INV_X1 port map( A => B(17), ZN => n48);
   U53 : INV_X1 port map( A => B(21), ZN => n44);
   U54 : INV_X1 port map( A => B(24), ZN => n41);
   U55 : INV_X1 port map( A => B(25), ZN => n40);
   U56 : INV_X1 port map( A => B(28), ZN => n37);
   U57 : INV_X1 port map( A => B(29), ZN => n36);
   U58 : INV_X1 port map( A => B(7), ZN => n58);
   U59 : INV_X1 port map( A => B(11), ZN => n54);
   U60 : INV_X1 port map( A => B(15), ZN => n50);
   U61 : INV_X1 port map( A => B(19), ZN => n46);
   U62 : INV_X1 port map( A => B(23), ZN => n42);
   U63 : INV_X1 port map( A => B(27), ZN => n38);
   U64 : INV_X1 port map( A => n159, ZN => GE_port);
   U65 : NAND2_X1 port map( A1 => GE_port, A2 => LE_port, ZN => NE);
   U66 : OAI21_X1 port map( B1 => n66, B2 => n67, A => n68, ZN => n65);
   U67 : MUX2_X1 port map( A => n69, B => n70, S => n3, Z => n68);
   U68 : NAND2_X1 port map( A1 => TC, A2 => B(31), ZN => n70);
   U69 : OR2_X1 port map( A1 => B(31), A2 => TC, ZN => n69);
   U70 : AOI22_X1 port map( A1 => A(30), A2 => n35, B1 => n71, B2 => n72, ZN =>
                           n66);
   U71 : AOI21_X1 port map( B1 => n73, B2 => n74, A => n75, ZN => n71);
   U72 : OAI211_X1 port map( C1 => n76, C2 => n77, A => n78, B => n79, ZN => 
                           n74);
   U73 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => n77);
   U74 : AOI211_X1 port map( C1 => n82, C2 => n83, A => n7, B => n84, ZN => n76
                           );
   U75 : OAI211_X1 port map( C1 => n86, C2 => n87, A => n88, B => n89, ZN => 
                           n83);
   U76 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => n87);
   U77 : AOI211_X1 port map( C1 => n92, C2 => n93, A => n11, B => n94, ZN => 
                           n86);
   U78 : OAI211_X1 port map( C1 => n96, C2 => n97, A => n98, B => n99, ZN => 
                           n93);
   U79 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => n97);
   U80 : AOI211_X1 port map( C1 => n102, C2 => n103, A => n15, B => n104, ZN =>
                           n96);
   U81 : OAI211_X1 port map( C1 => n106, C2 => n107, A => n108, B => n109, ZN 
                           => n103);
   U82 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => n107);
   U83 : AOI211_X1 port map( C1 => n112, C2 => n113, A => n19, B => n114, ZN =>
                           n106);
   U84 : OAI211_X1 port map( C1 => n116, C2 => n117, A => n118, B => n119, ZN 
                           => n113);
   U85 : NAND2_X1 port map( A1 => n120, A2 => n121, ZN => n117);
   U86 : AOI211_X1 port map( C1 => n122, C2 => n123, A => n23, B => n124, ZN =>
                           n116);
   U87 : OAI211_X1 port map( C1 => n126, C2 => n127, A => n128, B => n129, ZN 
                           => n123);
   U88 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => n127);
   U89 : AOI211_X1 port map( C1 => n132, C2 => n133, A => n27, B => n134, ZN =>
                           n126);
   U90 : NAND3_X1 port map( A1 => n136, A2 => n137, A3 => n138, ZN => n133);
   U91 : NAND3_X1 port map( A1 => n139, A2 => n140, A3 => n141, ZN => n136);
   U92 : OAI211_X1 port map( C1 => A(1), C2 => n34, A => n142, B => n143, ZN =>
                           n141);
   U93 : OAI21_X1 port map( B1 => n33, B2 => n144, A => B(1), ZN => n142);
   U94 : NAND2_X1 port map( A1 => A(0), A2 => n64, ZN => n144);
   U95 : NOR2_X1 port map( A1 => n145, A2 => n146, ZN => n132);
   U96 : NOR2_X1 port map( A1 => n147, A2 => n148, ZN => n122);
   U97 : NOR2_X1 port map( A1 => n149, A2 => n150, ZN => n112);
   U98 : NOR2_X1 port map( A1 => n151, A2 => n152, ZN => n102);
   U99 : NOR2_X1 port map( A1 => n153, A2 => n154, ZN => n92);
   U100 : NOR2_X1 port map( A1 => n155, A2 => n156, ZN => n82);
   U101 : NOR2_X1 port map( A1 => n157, A2 => n158, ZN => n73);
   U102 : OAI21_X1 port map( B1 => n160, B2 => n67, A => n161, ZN => n159);
   U103 : MUX2_X1 port map( A => n162, B => n163, S => TC, Z => n161);
   U104 : OR2_X1 port map( A1 => n3, A2 => B(31), ZN => n163);
   U105 : NAND2_X1 port map( A1 => B(31), A2 => n3, ZN => n162);
   U106 : XNOR2_X1 port map( A => n3, B => B(31), ZN => n67);
   U107 : AOI22_X1 port map( A1 => B(30), A2 => n4, B1 => n164, B2 => n72, ZN 
                           => n160);
   U108 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n72);
   U109 : AOI21_X1 port map( B1 => n165, B2 => n5, A => n158, ZN => n164);
   U110 : AND2_X1 port map( A1 => A(29), A2 => n36, ZN => n158);
   U111 : NOR2_X1 port map( A1 => n36, A2 => A(29), ZN => n75);
   U112 : AOI21_X1 port map( B1 => n166, B2 => n79, A => n167, ZN => n165);
   U113 : NOR2_X1 port map( A1 => n167, A2 => n157, ZN => n79);
   U114 : AND2_X1 port map( A1 => A(28), A2 => n37, ZN => n157);
   U115 : NOR2_X1 port map( A1 => n37, A2 => A(28), ZN => n167);
   U116 : AOI21_X1 port map( B1 => n168, B2 => n78, A => n6, ZN => n166);
   U117 : NAND2_X1 port map( A1 => A(27), A2 => n38, ZN => n80);
   U118 : OR2_X1 port map( A1 => n38, A2 => A(27), ZN => n78);
   U119 : AOI21_X1 port map( B1 => n169, B2 => n85, A => n170, ZN => n168);
   U120 : NOR2_X1 port map( A1 => n170, A2 => n8, ZN => n85);
   U121 : NAND2_X1 port map( A1 => A(26), A2 => n39, ZN => n81);
   U122 : NOR2_X1 port map( A1 => n39, A2 => A(26), ZN => n170);
   U123 : AOI21_X1 port map( B1 => n171, B2 => n9, A => n156, ZN => n169);
   U124 : AND2_X1 port map( A1 => A(25), A2 => n40, ZN => n156);
   U125 : NOR2_X1 port map( A1 => n40, A2 => A(25), ZN => n84);
   U126 : AOI21_X1 port map( B1 => n172, B2 => n89, A => n173, ZN => n171);
   U127 : NOR2_X1 port map( A1 => n173, A2 => n155, ZN => n89);
   U128 : AND2_X1 port map( A1 => A(24), A2 => n41, ZN => n155);
   U129 : NOR2_X1 port map( A1 => n41, A2 => A(24), ZN => n173);
   U130 : AOI21_X1 port map( B1 => n174, B2 => n88, A => n10, ZN => n172);
   U131 : NAND2_X1 port map( A1 => A(23), A2 => n42, ZN => n90);
   U132 : OR2_X1 port map( A1 => n42, A2 => A(23), ZN => n88);
   U133 : AOI21_X1 port map( B1 => n175, B2 => n95, A => n176, ZN => n174);
   U134 : NOR2_X1 port map( A1 => n176, A2 => n12, ZN => n95);
   U135 : NAND2_X1 port map( A1 => A(22), A2 => n43, ZN => n91);
   U136 : NOR2_X1 port map( A1 => n43, A2 => A(22), ZN => n176);
   U137 : AOI21_X1 port map( B1 => n177, B2 => n13, A => n154, ZN => n175);
   U138 : AND2_X1 port map( A1 => A(21), A2 => n44, ZN => n154);
   U139 : NOR2_X1 port map( A1 => n44, A2 => A(21), ZN => n94);
   U140 : AOI21_X1 port map( B1 => n178, B2 => n99, A => n179, ZN => n177);
   U141 : NOR2_X1 port map( A1 => n179, A2 => n153, ZN => n99);
   U142 : AND2_X1 port map( A1 => A(20), A2 => n45, ZN => n153);
   U143 : NOR2_X1 port map( A1 => n45, A2 => A(20), ZN => n179);
   U144 : AOI21_X1 port map( B1 => n180, B2 => n98, A => n14, ZN => n178);
   U145 : NAND2_X1 port map( A1 => A(19), A2 => n46, ZN => n100);
   U146 : OR2_X1 port map( A1 => n46, A2 => A(19), ZN => n98);
   U147 : AOI21_X1 port map( B1 => n181, B2 => n105, A => n182, ZN => n180);
   U148 : NOR2_X1 port map( A1 => n182, A2 => n16, ZN => n105);
   U149 : NAND2_X1 port map( A1 => A(18), A2 => n47, ZN => n101);
   U150 : NOR2_X1 port map( A1 => n47, A2 => A(18), ZN => n182);
   U151 : AOI21_X1 port map( B1 => n183, B2 => n17, A => n152, ZN => n181);
   U152 : AND2_X1 port map( A1 => A(17), A2 => n48, ZN => n152);
   U153 : NOR2_X1 port map( A1 => n48, A2 => A(17), ZN => n104);
   U154 : AOI21_X1 port map( B1 => n184, B2 => n109, A => n185, ZN => n183);
   U155 : NOR2_X1 port map( A1 => n185, A2 => n151, ZN => n109);
   U156 : AND2_X1 port map( A1 => A(16), A2 => n49, ZN => n151);
   U157 : NOR2_X1 port map( A1 => n49, A2 => A(16), ZN => n185);
   U158 : AOI21_X1 port map( B1 => n186, B2 => n108, A => n18, ZN => n184);
   U159 : NAND2_X1 port map( A1 => A(15), A2 => n50, ZN => n110);
   U160 : OR2_X1 port map( A1 => n50, A2 => A(15), ZN => n108);
   U161 : AOI21_X1 port map( B1 => n187, B2 => n115, A => n188, ZN => n186);
   U162 : NOR2_X1 port map( A1 => n188, A2 => n20, ZN => n115);
   U163 : NAND2_X1 port map( A1 => A(14), A2 => n51, ZN => n111);
   U164 : NOR2_X1 port map( A1 => n51, A2 => A(14), ZN => n188);
   U165 : AOI21_X1 port map( B1 => n189, B2 => n21, A => n150, ZN => n187);
   U166 : AND2_X1 port map( A1 => A(13), A2 => n52, ZN => n150);
   U167 : NOR2_X1 port map( A1 => n52, A2 => A(13), ZN => n114);
   U168 : AOI21_X1 port map( B1 => n190, B2 => n119, A => n191, ZN => n189);
   U169 : NOR2_X1 port map( A1 => n191, A2 => n149, ZN => n119);
   U170 : AND2_X1 port map( A1 => A(12), A2 => n53, ZN => n149);
   U171 : NOR2_X1 port map( A1 => n53, A2 => A(12), ZN => n191);
   U172 : AOI21_X1 port map( B1 => n192, B2 => n118, A => n22, ZN => n190);
   U173 : NAND2_X1 port map( A1 => A(11), A2 => n54, ZN => n120);
   U174 : OR2_X1 port map( A1 => n54, A2 => A(11), ZN => n118);
   U175 : AOI21_X1 port map( B1 => n193, B2 => n125, A => n194, ZN => n192);
   U176 : NOR2_X1 port map( A1 => n194, A2 => n24, ZN => n125);
   U177 : NAND2_X1 port map( A1 => A(10), A2 => n55, ZN => n121);
   U178 : NOR2_X1 port map( A1 => n55, A2 => A(10), ZN => n194);
   U179 : AOI21_X1 port map( B1 => n195, B2 => n25, A => n148, ZN => n193);
   U180 : AND2_X1 port map( A1 => A(9), A2 => n56, ZN => n148);
   U181 : NOR2_X1 port map( A1 => n56, A2 => A(9), ZN => n124);
   U182 : AOI21_X1 port map( B1 => n196, B2 => n129, A => n197, ZN => n195);
   U183 : NOR2_X1 port map( A1 => n197, A2 => n147, ZN => n129);
   U184 : AND2_X1 port map( A1 => A(8), A2 => n57, ZN => n147);
   U185 : NOR2_X1 port map( A1 => n57, A2 => A(8), ZN => n197);
   U186 : AOI21_X1 port map( B1 => n198, B2 => n128, A => n26, ZN => n196);
   U187 : NAND2_X1 port map( A1 => A(7), A2 => n58, ZN => n130);
   U188 : OR2_X1 port map( A1 => n58, A2 => A(7), ZN => n128);
   U189 : AOI21_X1 port map( B1 => n199, B2 => n135, A => n200, ZN => n198);
   U190 : NOR2_X1 port map( A1 => n200, A2 => n28, ZN => n135);
   U191 : NAND2_X1 port map( A1 => A(6), A2 => n59, ZN => n131);
   U192 : NOR2_X1 port map( A1 => n59, A2 => A(6), ZN => n200);
   U193 : AOI21_X1 port map( B1 => n201, B2 => n29, A => n146, ZN => n199);
   U194 : AND2_X1 port map( A1 => A(5), A2 => n60, ZN => n146);
   U195 : NOR2_X1 port map( A1 => n60, A2 => A(5), ZN => n134);
   U196 : AOI21_X1 port map( B1 => n202, B2 => n138, A => n203, ZN => n201);
   U197 : NOR2_X1 port map( A1 => n203, A2 => n145, ZN => n138);
   U198 : AND2_X1 port map( A1 => A(4), A2 => n61, ZN => n145);
   U199 : NOR2_X1 port map( A1 => n61, A2 => A(4), ZN => n203);
   U200 : AOI21_X1 port map( B1 => n204, B2 => n137, A => n30, ZN => n202);
   U201 : NAND2_X1 port map( A1 => A(3), A2 => n62, ZN => n139);
   U202 : OR2_X1 port map( A1 => n62, A2 => A(3), ZN => n137);
   U203 : AOI21_X1 port map( B1 => n32, B2 => n143, A => n205, ZN => n204);
   U204 : NOR2_X1 port map( A1 => n205, A2 => n31, ZN => n143);
   U205 : NAND2_X1 port map( A1 => A(2), A2 => n63, ZN => n140);
   U206 : NOR2_X1 port map( A1 => n63, A2 => A(2), ZN => n205);
   U207 : OAI22_X1 port map( A1 => n207, A2 => B(1), B1 => n33, B2 => n208, ZN 
                           => n206);
   U208 : AND2_X1 port map( A1 => n208, A2 => n33, ZN => n207);
   U209 : NOR2_X1 port map( A1 => n64, A2 => A(0), ZN => n208);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_addsub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in std_logic;
         SUM : out std_logic_vector (31 downto 0);  CO : out std_logic);

end ALU_N32_DW01_addsub_0;

architecture SYN_rpl of ALU_N32_DW01_addsub_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, B_AS_31_port, 
      B_AS_30_port, B_AS_29_port, B_AS_28_port, B_AS_27_port, B_AS_26_port, 
      B_AS_25_port, B_AS_24_port, B_AS_23_port, B_AS_22_port, B_AS_21_port, 
      B_AS_20_port, B_AS_19_port, B_AS_18_port, B_AS_17_port, B_AS_16_port, 
      B_AS_15_port, B_AS_14_port, B_AS_13_port, B_AS_12_port, B_AS_11_port, 
      B_AS_10_port, B_AS_9_port, B_AS_8_port, B_AS_7_port, B_AS_6_port, 
      B_AS_5_port, B_AS_4_port, B_AS_3_port, B_AS_2_port, B_AS_1_port, 
      B_AS_0_port, n_1039 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B_AS_31_port, CI => carry_31_port, 
                           CO => n_1039, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B_AS_30_port, CI => carry_30_port, 
                           CO => carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B_AS_29_port, CI => carry_29_port, 
                           CO => carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B_AS_28_port, CI => carry_28_port, 
                           CO => carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B_AS_27_port, CI => carry_27_port, 
                           CO => carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B_AS_26_port, CI => carry_26_port, 
                           CO => carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B_AS_25_port, CI => carry_25_port, 
                           CO => carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B_AS_24_port, CI => carry_24_port, 
                           CO => carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B_AS_23_port, CI => carry_23_port, 
                           CO => carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B_AS_22_port, CI => carry_22_port, 
                           CO => carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B_AS_21_port, CI => carry_21_port, 
                           CO => carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B_AS_20_port, CI => carry_20_port, 
                           CO => carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B_AS_19_port, CI => carry_19_port, 
                           CO => carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B_AS_18_port, CI => carry_18_port, 
                           CO => carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B_AS_17_port, CI => carry_17_port, 
                           CO => carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B_AS_16_port, CI => carry_16_port, 
                           CO => carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B_AS_15_port, CI => carry_15_port, 
                           CO => carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B_AS_14_port, CI => carry_14_port, 
                           CO => carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B_AS_13_port, CI => carry_13_port, 
                           CO => carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B_AS_12_port, CI => carry_12_port, 
                           CO => carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B_AS_11_port, CI => carry_11_port, 
                           CO => carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B_AS_10_port, CI => carry_10_port, 
                           CO => carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B_AS_9_port, CI => carry_9_port, CO 
                           => carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B_AS_8_port, CI => carry_8_port, CO 
                           => carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B_AS_7_port, CI => carry_7_port, CO 
                           => carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B_AS_6_port, CI => carry_6_port, CO 
                           => carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B_AS_5_port, CI => carry_5_port, CO 
                           => carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B_AS_4_port, CI => carry_4_port, CO 
                           => carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B_AS_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B_AS_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B_AS_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_AS_9_port);
   U2 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_AS_8_port);
   U3 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_AS_7_port);
   U4 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_AS_6_port);
   U5 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_AS_5_port);
   U6 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_AS_4_port);
   U7 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_AS_3_port);
   U8 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_AS_31_port);
   U9 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_AS_30_port);
   U10 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_AS_2_port);
   U11 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_AS_29_port);
   U12 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_AS_28_port);
   U13 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_AS_27_port);
   U14 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_AS_26_port);
   U15 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_AS_25_port);
   U16 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_AS_24_port);
   U17 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_AS_23_port);
   U18 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_AS_22_port);
   U19 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_AS_21_port);
   U20 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_AS_20_port);
   U21 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_AS_1_port);
   U22 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_AS_19_port);
   U23 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_AS_18_port);
   U24 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_AS_17_port);
   U25 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_AS_16_port);
   U26 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_AS_15_port);
   U27 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_AS_14_port);
   U28 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_AS_13_port);
   U29 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_AS_12_port);
   U30 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_AS_11_port);
   U31 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_AS_10_port);
   U32 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_31 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_31;

architecture SYN_BEHAVIOUR of NAND4_31 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_30 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_30;

architecture SYN_BEHAVIOUR of NAND4_30 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_29 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_29;

architecture SYN_BEHAVIOUR of NAND4_29 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_28 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_28;

architecture SYN_BEHAVIOUR of NAND4_28 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_27 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_27;

architecture SYN_BEHAVIOUR of NAND4_27 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_26 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_26;

architecture SYN_BEHAVIOUR of NAND4_26 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_25 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_25;

architecture SYN_BEHAVIOUR of NAND4_25 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_24 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_24;

architecture SYN_BEHAVIOUR of NAND4_24 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_23 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_23;

architecture SYN_BEHAVIOUR of NAND4_23 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_22 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_22;

architecture SYN_BEHAVIOUR of NAND4_22 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_21 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_21;

architecture SYN_BEHAVIOUR of NAND4_21 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_20 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_20;

architecture SYN_BEHAVIOUR of NAND4_20 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_19 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_19;

architecture SYN_BEHAVIOUR of NAND4_19 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_18 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_18;

architecture SYN_BEHAVIOUR of NAND4_18 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_17 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_17;

architecture SYN_BEHAVIOUR of NAND4_17 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_16 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_16;

architecture SYN_BEHAVIOUR of NAND4_16 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_15 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_15;

architecture SYN_BEHAVIOUR of NAND4_15 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_14 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_14;

architecture SYN_BEHAVIOUR of NAND4_14 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_13 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_13;

architecture SYN_BEHAVIOUR of NAND4_13 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_12 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_12;

architecture SYN_BEHAVIOUR of NAND4_12 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_11 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_11;

architecture SYN_BEHAVIOUR of NAND4_11 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_10 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_10;

architecture SYN_BEHAVIOUR of NAND4_10 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_9 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_9;

architecture SYN_BEHAVIOUR of NAND4_9 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_8 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_8;

architecture SYN_BEHAVIOUR of NAND4_8 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_7 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_7;

architecture SYN_BEHAVIOUR of NAND4_7 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_6 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_6;

architecture SYN_BEHAVIOUR of NAND4_6 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_5 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_5;

architecture SYN_BEHAVIOUR of NAND4_5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_4 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_4;

architecture SYN_BEHAVIOUR of NAND4_4 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_3 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_3;

architecture SYN_BEHAVIOUR of NAND4_3 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_2 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_2;

architecture SYN_BEHAVIOUR of NAND4_2 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_1 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_1;

architecture SYN_BEHAVIOUR of NAND4_1 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_127 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_127;

architecture SYN_BEHAVIOUR of NAND3_127 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_126 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_126;

architecture SYN_BEHAVIOUR of NAND3_126 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_125 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_125;

architecture SYN_BEHAVIOUR of NAND3_125 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_124 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_124;

architecture SYN_BEHAVIOUR of NAND3_124 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_123 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_123;

architecture SYN_BEHAVIOUR of NAND3_123 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_122 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_122;

architecture SYN_BEHAVIOUR of NAND3_122 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_121 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_121;

architecture SYN_BEHAVIOUR of NAND3_121 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_120 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_120;

architecture SYN_BEHAVIOUR of NAND3_120 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_119 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_119;

architecture SYN_BEHAVIOUR of NAND3_119 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_118 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_118;

architecture SYN_BEHAVIOUR of NAND3_118 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_117 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_117;

architecture SYN_BEHAVIOUR of NAND3_117 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_116 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_116;

architecture SYN_BEHAVIOUR of NAND3_116 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_115 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_115;

architecture SYN_BEHAVIOUR of NAND3_115 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_114 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_114;

architecture SYN_BEHAVIOUR of NAND3_114 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_113 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_113;

architecture SYN_BEHAVIOUR of NAND3_113 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_112 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_112;

architecture SYN_BEHAVIOUR of NAND3_112 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_111 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_111;

architecture SYN_BEHAVIOUR of NAND3_111 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_110 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_110;

architecture SYN_BEHAVIOUR of NAND3_110 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_109 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_109;

architecture SYN_BEHAVIOUR of NAND3_109 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_108 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_108;

architecture SYN_BEHAVIOUR of NAND3_108 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_107 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_107;

architecture SYN_BEHAVIOUR of NAND3_107 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_106 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_106;

architecture SYN_BEHAVIOUR of NAND3_106 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_105 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_105;

architecture SYN_BEHAVIOUR of NAND3_105 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_104 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_104;

architecture SYN_BEHAVIOUR of NAND3_104 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_103 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_103;

architecture SYN_BEHAVIOUR of NAND3_103 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_102 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_102;

architecture SYN_BEHAVIOUR of NAND3_102 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_101 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_101;

architecture SYN_BEHAVIOUR of NAND3_101 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_100 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_100;

architecture SYN_BEHAVIOUR of NAND3_100 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_99 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_99;

architecture SYN_BEHAVIOUR of NAND3_99 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_98 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_98;

architecture SYN_BEHAVIOUR of NAND3_98 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_97 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_97;

architecture SYN_BEHAVIOUR of NAND3_97 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_96 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_96;

architecture SYN_BEHAVIOUR of NAND3_96 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_95 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_95;

architecture SYN_BEHAVIOUR of NAND3_95 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_94 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_94;

architecture SYN_BEHAVIOUR of NAND3_94 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_93 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_93;

architecture SYN_BEHAVIOUR of NAND3_93 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_92 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_92;

architecture SYN_BEHAVIOUR of NAND3_92 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_91 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_91;

architecture SYN_BEHAVIOUR of NAND3_91 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_90 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_90;

architecture SYN_BEHAVIOUR of NAND3_90 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_89 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_89;

architecture SYN_BEHAVIOUR of NAND3_89 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_88 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_88;

architecture SYN_BEHAVIOUR of NAND3_88 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_87 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_87;

architecture SYN_BEHAVIOUR of NAND3_87 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_86 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_86;

architecture SYN_BEHAVIOUR of NAND3_86 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_85 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_85;

architecture SYN_BEHAVIOUR of NAND3_85 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_84 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_84;

architecture SYN_BEHAVIOUR of NAND3_84 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_83 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_83;

architecture SYN_BEHAVIOUR of NAND3_83 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_82 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_82;

architecture SYN_BEHAVIOUR of NAND3_82 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_81 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_81;

architecture SYN_BEHAVIOUR of NAND3_81 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_80 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_80;

architecture SYN_BEHAVIOUR of NAND3_80 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_79 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_79;

architecture SYN_BEHAVIOUR of NAND3_79 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_78 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_78;

architecture SYN_BEHAVIOUR of NAND3_78 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_77 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_77;

architecture SYN_BEHAVIOUR of NAND3_77 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_76 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_76;

architecture SYN_BEHAVIOUR of NAND3_76 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_75 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_75;

architecture SYN_BEHAVIOUR of NAND3_75 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_74 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_74;

architecture SYN_BEHAVIOUR of NAND3_74 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_73 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_73;

architecture SYN_BEHAVIOUR of NAND3_73 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_72 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_72;

architecture SYN_BEHAVIOUR of NAND3_72 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_71 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_71;

architecture SYN_BEHAVIOUR of NAND3_71 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_70 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_70;

architecture SYN_BEHAVIOUR of NAND3_70 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_69 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_69;

architecture SYN_BEHAVIOUR of NAND3_69 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_68 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_68;

architecture SYN_BEHAVIOUR of NAND3_68 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_67 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_67;

architecture SYN_BEHAVIOUR of NAND3_67 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_66 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_66;

architecture SYN_BEHAVIOUR of NAND3_66 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_65 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_65;

architecture SYN_BEHAVIOUR of NAND3_65 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_64 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_64;

architecture SYN_BEHAVIOUR of NAND3_64 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_63 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_63;

architecture SYN_BEHAVIOUR of NAND3_63 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_62 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_62;

architecture SYN_BEHAVIOUR of NAND3_62 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_61 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_61;

architecture SYN_BEHAVIOUR of NAND3_61 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_60 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_60;

architecture SYN_BEHAVIOUR of NAND3_60 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_59 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_59;

architecture SYN_BEHAVIOUR of NAND3_59 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_58 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_58;

architecture SYN_BEHAVIOUR of NAND3_58 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_57 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_57;

architecture SYN_BEHAVIOUR of NAND3_57 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_56 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_56;

architecture SYN_BEHAVIOUR of NAND3_56 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_55 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_55;

architecture SYN_BEHAVIOUR of NAND3_55 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_54 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_54;

architecture SYN_BEHAVIOUR of NAND3_54 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_53 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_53;

architecture SYN_BEHAVIOUR of NAND3_53 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_52 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_52;

architecture SYN_BEHAVIOUR of NAND3_52 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_51 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_51;

architecture SYN_BEHAVIOUR of NAND3_51 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_50 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_50;

architecture SYN_BEHAVIOUR of NAND3_50 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_49 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_49;

architecture SYN_BEHAVIOUR of NAND3_49 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_48 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_48;

architecture SYN_BEHAVIOUR of NAND3_48 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_47 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_47;

architecture SYN_BEHAVIOUR of NAND3_47 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_46 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_46;

architecture SYN_BEHAVIOUR of NAND3_46 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_45 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_45;

architecture SYN_BEHAVIOUR of NAND3_45 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_44 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_44;

architecture SYN_BEHAVIOUR of NAND3_44 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_43 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_43;

architecture SYN_BEHAVIOUR of NAND3_43 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_42 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_42;

architecture SYN_BEHAVIOUR of NAND3_42 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_41 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_41;

architecture SYN_BEHAVIOUR of NAND3_41 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_40 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_40;

architecture SYN_BEHAVIOUR of NAND3_40 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_39 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_39;

architecture SYN_BEHAVIOUR of NAND3_39 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_38 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_38;

architecture SYN_BEHAVIOUR of NAND3_38 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_37 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_37;

architecture SYN_BEHAVIOUR of NAND3_37 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_36 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_36;

architecture SYN_BEHAVIOUR of NAND3_36 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_35 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_35;

architecture SYN_BEHAVIOUR of NAND3_35 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_34 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_34;

architecture SYN_BEHAVIOUR of NAND3_34 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_33 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_33;

architecture SYN_BEHAVIOUR of NAND3_33 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_32 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_32;

architecture SYN_BEHAVIOUR of NAND3_32 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_31 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_31;

architecture SYN_BEHAVIOUR of NAND3_31 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_30 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_30;

architecture SYN_BEHAVIOUR of NAND3_30 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_29 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_29;

architecture SYN_BEHAVIOUR of NAND3_29 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_28 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_28;

architecture SYN_BEHAVIOUR of NAND3_28 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_27 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_27;

architecture SYN_BEHAVIOUR of NAND3_27 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_26 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_26;

architecture SYN_BEHAVIOUR of NAND3_26 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_25 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_25;

architecture SYN_BEHAVIOUR of NAND3_25 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_24 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_24;

architecture SYN_BEHAVIOUR of NAND3_24 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_23 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_23;

architecture SYN_BEHAVIOUR of NAND3_23 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_22 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_22;

architecture SYN_BEHAVIOUR of NAND3_22 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_21 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_21;

architecture SYN_BEHAVIOUR of NAND3_21 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_20 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_20;

architecture SYN_BEHAVIOUR of NAND3_20 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_19 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_19;

architecture SYN_BEHAVIOUR of NAND3_19 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_18 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_18;

architecture SYN_BEHAVIOUR of NAND3_18 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_17 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_17;

architecture SYN_BEHAVIOUR of NAND3_17 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_16 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_16;

architecture SYN_BEHAVIOUR of NAND3_16 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_15 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_15;

architecture SYN_BEHAVIOUR of NAND3_15 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_14 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_14;

architecture SYN_BEHAVIOUR of NAND3_14 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_13 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_13;

architecture SYN_BEHAVIOUR of NAND3_13 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_12 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_12;

architecture SYN_BEHAVIOUR of NAND3_12 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_11 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_11;

architecture SYN_BEHAVIOUR of NAND3_11 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_10 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_10;

architecture SYN_BEHAVIOUR of NAND3_10 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_9 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_9;

architecture SYN_BEHAVIOUR of NAND3_9 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_8 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_8;

architecture SYN_BEHAVIOUR of NAND3_8 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_7 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_7;

architecture SYN_BEHAVIOUR of NAND3_7 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_6 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_6;

architecture SYN_BEHAVIOUR of NAND3_6 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_5 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_5;

architecture SYN_BEHAVIOUR of NAND3_5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_4 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_4;

architecture SYN_BEHAVIOUR of NAND3_4 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_3 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_3;

architecture SYN_BEHAVIOUR of NAND3_3 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_2 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_2;

architecture SYN_BEHAVIOUR of NAND3_2 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_1 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_1;

architecture SYN_BEHAVIOUR of NAND3_1 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT5_1 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_GENERIC_NBIT5_1;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT5_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U5 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_4;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_3;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n33, n34, n35 : std_logic;

begin
   
   U1 : BUF_X4 port map( A => n35, Z => Y(0));
   U2 : BUF_X4 port map( A => n34, Z => Y(1));
   U3 : BUF_X4 port map( A => n33, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U5 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U6 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U7 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U8 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U9 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U10 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U11 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U12 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U13 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U14 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U15 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U16 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U17 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U20 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U23 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U24 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U25 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U26 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U27 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U28 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U29 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U30 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U31 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U32 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U33 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => n33);
   U34 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => n34);
   U35 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_2;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_1;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT5_2 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 downto 
         0);  DATA_OUT : out std_logic_vector (4 downto 0));

end REG_GENERIC_NBIT5_2;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT5_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n14, CK => CLK, Q => DATA_OUT(4)
                           , QN => n13);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n15, CK => CLK, Q => DATA_OUT(3)
                           , QN => n12);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n16, CK => CLK, Q => DATA_OUT(2)
                           , QN => n11);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n17, CK => CLK, Q => DATA_OUT(1)
                           , QN => n10);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n18, CK => CLK, Q => DATA_OUT(0)
                           , QN => n9);
   U3 : OAI21_X1 port map( B1 => n13, B2 => n1, A => n2, ZN => n14);
   U4 : NAND2_X1 port map( A1 => DATA_IN(4), A2 => n3, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n12, B2 => n1, A => n4, ZN => n15);
   U6 : NAND2_X1 port map( A1 => DATA_IN(3), A2 => n3, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n11, B2 => n1, A => n5, ZN => n16);
   U8 : NAND2_X1 port map( A1 => DATA_IN(2), A2 => n3, ZN => n5);
   U9 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n6, ZN => n17);
   U10 : NAND2_X1 port map( A1 => DATA_IN(1), A2 => n3, ZN => n6);
   U11 : OAI21_X1 port map( B1 => n9, B2 => n1, A => n7, ZN => n18);
   U12 : NAND2_X1 port map( A1 => DATA_IN(0), A2 => n3, ZN => n7);
   U13 : AND2_X1 port map( A1 => RST, A2 => n1, ZN => n3);
   U14 : NAND2_X1 port map( A1 => n8, A2 => RST, ZN => n1);
   U15 : INV_X1 port map( A => EN, ZN => n8);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT5_1 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 downto 
         0);  DATA_OUT : out std_logic_vector (4 downto 0));

end REG_GENERIC_NBIT5_1;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n14, CK => CLK, Q => DATA_OUT(4)
                           , QN => n13);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n15, CK => CLK, Q => DATA_OUT(3)
                           , QN => n12);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n16, CK => CLK, Q => DATA_OUT(2)
                           , QN => n11);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n17, CK => CLK, Q => DATA_OUT(1)
                           , QN => n10);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n18, CK => CLK, Q => DATA_OUT(0)
                           , QN => n9);
   U3 : OAI21_X1 port map( B1 => n13, B2 => n1, A => n2, ZN => n14);
   U4 : NAND2_X1 port map( A1 => DATA_IN(4), A2 => n3, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n12, B2 => n1, A => n4, ZN => n15);
   U6 : NAND2_X1 port map( A1 => DATA_IN(3), A2 => n3, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n11, B2 => n1, A => n5, ZN => n16);
   U8 : NAND2_X1 port map( A1 => DATA_IN(2), A2 => n3, ZN => n5);
   U9 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n6, ZN => n17);
   U10 : NAND2_X1 port map( A1 => DATA_IN(1), A2 => n3, ZN => n6);
   U11 : OAI21_X1 port map( B1 => n9, B2 => n1, A => n7, ZN => n18);
   U12 : NAND2_X1 port map( A1 => DATA_IN(0), A2 => n3, ZN => n7);
   U13 : AND2_X1 port map( A1 => RST, A2 => n1, ZN => n3);
   U14 : NAND2_X1 port map( A1 => n8, A2 => RST, ZN => n1);
   U15 : INV_X1 port map( A => EN, ZN => n8);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_8 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_8;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_7 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_7;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_6 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_6;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_5 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_5;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_4 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_4;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045
      , n_1046, n_1047, n_1048, n_1049 : std_logic;

begin
   DATA_OUT <= ( DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port );
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n60, CK => CLK, Q => 
                           DATA_OUT_31_port, QN => n59);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n61, CK => CLK, Q => 
                           DATA_OUT_30_port, QN => n58);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n62, CK => CLK, Q => 
                           DATA_OUT_29_port, QN => n57);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n63, CK => CLK, Q => 
                           DATA_OUT_28_port, QN => n56);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n64, CK => CLK, Q => 
                           DATA_OUT_27_port, QN => n55);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n65, CK => CLK, Q => 
                           DATA_OUT_26_port, QN => n54);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n66, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_1040);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n67, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n_1041);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_1042);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n_1043);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n_1044);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_1045);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_1046);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_1047);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_1048);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n_1049);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n53);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n52);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n51);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n50);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n49);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n48);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n47);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n46);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n45);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n44);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT_5_port, QN => n43);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n42);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n41);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n40);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n90, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n39);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n91, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n38);
   U3 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n3, ZN => n60);
   U4 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U5 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n4, ZN => n61);
   U6 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U7 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n5, ZN => n62);
   U8 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U9 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n6, ZN => n63);
   U10 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U11 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n7, ZN => n64)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U13 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n8, ZN => n65)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U15 : INV_X1 port map( A => n9, ZN => n66);
   U16 : AOI22_X1 port map( A1 => DATA_IN(25), A2 => n10, B1 => 
                           DATA_OUT_25_port, B2 => n11, ZN => n9);
   U17 : INV_X1 port map( A => n12, ZN => n67);
   U18 : AOI22_X1 port map( A1 => DATA_IN(24), A2 => n10, B1 => 
                           DATA_OUT_24_port, B2 => n11, ZN => n12);
   U19 : INV_X1 port map( A => n13, ZN => n68);
   U20 : AOI22_X1 port map( A1 => DATA_IN(23), A2 => n10, B1 => 
                           DATA_OUT_23_port, B2 => n11, ZN => n13);
   U21 : INV_X1 port map( A => n14, ZN => n69);
   U22 : AOI22_X1 port map( A1 => DATA_IN(22), A2 => n10, B1 => 
                           DATA_OUT_22_port, B2 => n11, ZN => n14);
   U23 : INV_X1 port map( A => n15, ZN => n70);
   U24 : AOI22_X1 port map( A1 => DATA_IN(21), A2 => n10, B1 => 
                           DATA_OUT_21_port, B2 => n11, ZN => n15);
   U25 : INV_X1 port map( A => n16, ZN => n71);
   U26 : AOI22_X1 port map( A1 => DATA_IN(20), A2 => n10, B1 => 
                           DATA_OUT_20_port, B2 => n11, ZN => n16);
   U27 : INV_X1 port map( A => n17, ZN => n72);
   U28 : AOI22_X1 port map( A1 => DATA_IN(19), A2 => n10, B1 => 
                           DATA_OUT_19_port, B2 => n11, ZN => n17);
   U29 : INV_X1 port map( A => n18, ZN => n73);
   U30 : AOI22_X1 port map( A1 => DATA_IN(18), A2 => n10, B1 => 
                           DATA_OUT_18_port, B2 => n11, ZN => n18);
   U31 : INV_X1 port map( A => n19, ZN => n74);
   U32 : AOI22_X1 port map( A1 => DATA_IN(17), A2 => n10, B1 => 
                           DATA_OUT_17_port, B2 => n11, ZN => n19);
   U33 : INV_X1 port map( A => n20, ZN => n75);
   U34 : AOI22_X1 port map( A1 => DATA_IN(16), A2 => n10, B1 => 
                           DATA_OUT_16_port, B2 => n11, ZN => n20);
   U35 : INV_X1 port map( A => n1, ZN => n11);
   U36 : INV_X1 port map( A => n2, ZN => n10);
   U37 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n21, ZN => n76
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n21);
   U39 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n22, ZN => n77
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n22);
   U41 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n23, ZN => n78
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n23);
   U43 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n24, ZN => n79
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n24);
   U45 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n25, ZN => n80
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n25);
   U47 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n26, ZN => n81
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n26);
   U49 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n27, ZN => n82
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n27);
   U51 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n28, ZN => n83
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n28);
   U53 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n29, ZN => n84
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n29);
   U55 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n30, ZN => n85
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n30);
   U57 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n31, ZN => n86
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n31);
   U59 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n32, ZN => n87
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n32);
   U61 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n33, ZN => n88
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n33);
   U63 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n34, ZN => n89
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n34);
   U65 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n35, ZN => n90
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n35);
   U67 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n36, ZN => n91
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n36);
   U69 : NAND2_X1 port map( A1 => RST, A2 => n1, ZN => n2);
   U70 : NAND2_X1 port map( A1 => n37, A2 => RST, ZN => n1);
   U71 : INV_X1 port map( A => EN, ZN => n37);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_3 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_3;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n90, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n91, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n92, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n93, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n83, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n84, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n85, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n68, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(0), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(31), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(30), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(29), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(28), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(27), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(26), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(25), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(24), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(23), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(14), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(13), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(12), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(11), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(10), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(9), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(8), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(7), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(15), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(22), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(21), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(20), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(19), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(18), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(17), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(16), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(6), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(5), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(4), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(3), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(2), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(1), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_2 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_2;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_1 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_1;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BARREL_SHIFTER_N32 is

   port( CONF : in std_logic;  DATA1, DATA2 : in std_logic_vector (31 downto 0)
         ;  OUTPUT : out std_logic_vector (31 downto 0));

end BARREL_SHIFTER_N32;

architecture SYN_BEHAVIOR of BARREL_SHIFTER_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal COARSE_39_port, COARSE_38_port, COARSE_37_port, COARSE_36_port, 
      COARSE_35_port, COARSE_34_port, COARSE_33_port, COARSE_32_port, 
      COARSE_31_port, COARSE_30_port, COARSE_29_port, COARSE_28_port, 
      COARSE_27_port, COARSE_26_port, COARSE_25_port, COARSE_24_port, 
      COARSE_23_port, COARSE_22_port, COARSE_21_port, COARSE_20_port, 
      COARSE_19_port, COARSE_18_port, COARSE_17_port, COARSE_16_port, 
      COARSE_15_port, COARSE_14_port, COARSE_13_port, COARSE_12_port, 
      COARSE_11_port, COARSE_10_port, COARSE_9_port, COARSE_8_port, 
      COARSE_7_port, COARSE_6_port, COARSE_5_port, COARSE_4_port, COARSE_3_port
      , COARSE_2_port, COARSE_1_port, COARSE_0_port, SL_OUT_31_port, 
      SL_OUT_30_port, SL_OUT_29_port, SL_OUT_28_port, SL_OUT_27_port, 
      SL_OUT_26_port, SL_OUT_25_port, SL_OUT_24_port, SL_OUT_23_port, 
      SL_OUT_22_port, SL_OUT_21_port, SL_OUT_20_port, SL_OUT_19_port, 
      SL_OUT_18_port, SL_OUT_17_port, SL_OUT_16_port, SL_OUT_15_port, 
      SL_OUT_14_port, SL_OUT_13_port, SL_OUT_12_port, SL_OUT_11_port, 
      SL_OUT_10_port, SL_OUT_9_port, SL_OUT_8_port, SL_OUT_7_port, 
      SL_OUT_6_port, SL_OUT_5_port, SL_OUT_4_port, SL_OUT_3_port, SL_OUT_2_port
      , SL_OUT_1_port, SL_OUT_0_port, SR_OUT_31_port, SR_OUT_30_port, 
      SR_OUT_29_port, SR_OUT_28_port, SR_OUT_27_port, SR_OUT_26_port, 
      SR_OUT_25_port, SR_OUT_24_port, SR_OUT_23_port, SR_OUT_22_port, 
      SR_OUT_21_port, SR_OUT_20_port, SR_OUT_19_port, SR_OUT_18_port, 
      SR_OUT_17_port, SR_OUT_16_port, SR_OUT_15_port, SR_OUT_14_port, 
      SR_OUT_13_port, SR_OUT_12_port, SR_OUT_11_port, SR_OUT_10_port, 
      SR_OUT_9_port, SR_OUT_8_port, SR_OUT_7_port, SR_OUT_6_port, SR_OUT_5_port
      , SR_OUT_4_port, SR_OUT_3_port, SR_OUT_2_port, SR_OUT_1_port, 
      SR_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325 : std_logic;

begin
   
   U2 : NOR3_X2 port map( A1 => n294, A2 => n241, A3 => n295, ZN => n255);
   U3 : NOR3_X4 port map( A1 => n241, A2 => DATA2(3), A3 => n294, ZN => n248);
   U4 : NOR3_X2 port map( A1 => n294, A2 => CONF, A3 => n295, ZN => n273);
   U5 : NAND3_X2 port map( A1 => n295, A2 => n294, A3 => CONF, ZN => n242);
   U6 : INV_X2 port map( A => CONF, ZN => n241);
   U7 : NOR3_X4 port map( A1 => CONF, A2 => DATA2(3), A3 => n294, ZN => n274);
   U8 : NOR3_X4 port map( A1 => CONF, A2 => DATA2(4), A3 => n295, ZN => n296);
   U9 : NOR3_X4 port map( A1 => DATA2(3), A2 => DATA2(4), A3 => CONF, ZN => 
                           n247);
   U10 : INV_X1 port map( A => COARSE_5_port, ZN => n162);
   U11 : INV_X1 port map( A => COARSE_4_port, ZN => n156);
   U12 : INV_X1 port map( A => COARSE_34_port, ZN => n146);
   U13 : INV_X1 port map( A => COARSE_35_port, ZN => n152);
   U14 : INV_X1 port map( A => n133, ZN => n164);
   U15 : INV_X1 port map( A => n12, ZN => n170);
   U16 : INV_X1 port map( A => n73, ZN => n211);
   U17 : INV_X1 port map( A => n69, ZN => n158);
   U18 : INV_X1 port map( A => COARSE_25_port, ZN => n145);
   U19 : INV_X1 port map( A => COARSE_24_port, ZN => n140);
   U20 : INV_X1 port map( A => COARSE_26_port, ZN => n150);
   U21 : INV_X1 port map( A => COARSE_27_port, ZN => n155);
   U22 : INV_X1 port map( A => COARSE_28_port, ZN => n161);
   U23 : INV_X1 port map( A => COARSE_29_port, ZN => n167);
   U24 : INV_X1 port map( A => COARSE_30_port, ZN => n196);
   U25 : INV_X1 port map( A => COARSE_31_port, ZN => n232);
   U26 : INV_X1 port map( A => COARSE_6_port, ZN => n168);
   U27 : INV_X1 port map( A => COARSE_7_port, ZN => n205);
   U28 : INV_X1 port map( A => COARSE_8_port, ZN => n137);
   U29 : INV_X1 port map( A => COARSE_9_port, ZN => n141);
   U30 : INV_X1 port map( A => COARSE_10_port, ZN => n149);
   U31 : INV_X1 port map( A => COARSE_11_port, ZN => n154);
   U32 : INV_X1 port map( A => COARSE_12_port, ZN => n160);
   U33 : INV_X1 port map( A => COARSE_13_port, ZN => n166);
   U34 : INV_X1 port map( A => COARSE_14_port, ZN => n187);
   U35 : INV_X1 port map( A => COARSE_15_port, ZN => n223);
   U36 : INV_X1 port map( A => COARSE_16_port, ZN => n139);
   U37 : INV_X1 port map( A => COARSE_17_port, ZN => n144);
   U38 : INV_X1 port map( A => COARSE_18_port, ZN => n148);
   U39 : INV_X1 port map( A => COARSE_19_port, ZN => n153);
   U40 : INV_X1 port map( A => COARSE_20_port, ZN => n159);
   U41 : INV_X1 port map( A => COARSE_21_port, ZN => n165);
   U42 : INV_X1 port map( A => COARSE_22_port, ZN => n178);
   U43 : INV_X1 port map( A => COARSE_23_port, ZN => n214);
   U44 : INV_X1 port map( A => COARSE_2_port, ZN => n147);
   U45 : INV_X1 port map( A => COARSE_3_port, ZN => n151);
   U46 : INV_X1 port map( A => COARSE_33_port, ZN => n142);
   U47 : INV_X1 port map( A => COARSE_32_port, ZN => n138);
   U48 : INV_X1 port map( A => COARSE_37_port, ZN => n163);
   U49 : INV_X1 port map( A => COARSE_36_port, ZN => n157);
   U50 : INV_X1 port map( A => n11, ZN => n206);
   U51 : INV_X1 port map( A => COARSE_1_port, ZN => n143);
   U52 : INV_X1 port map( A => n76, ZN => n173);
   U53 : INV_X1 port map( A => n14, ZN => n169);
   U54 : INV_X1 port map( A => n78, ZN => n210);
   U55 : INV_X1 port map( A => n16, ZN => n207);
   U56 : INV_X1 port map( A => n80, ZN => n174);
   U57 : INV_X1 port map( A => n18, ZN => n171);
   U58 : INV_X1 port map( A => n82, ZN => n212);
   U59 : INV_X1 port map( A => n20, ZN => n208);
   U60 : INV_X1 port map( A => n84, ZN => n175);
   U61 : INV_X1 port map( A => n22, ZN => n172);
   U62 : INV_X1 port map( A => n86, ZN => n213);
   U63 : INV_X1 port map( A => n24, ZN => n209);
   U64 : INV_X1 port map( A => n88, ZN => n192);
   U65 : INV_X1 port map( A => n26, ZN => n188);
   U66 : INV_X1 port map( A => n90, ZN => n228);
   U67 : INV_X1 port map( A => n28, ZN => n224);
   U68 : INV_X1 port map( A => n92, ZN => n193);
   U69 : INV_X1 port map( A => n30, ZN => n189);
   U70 : INV_X1 port map( A => n94, ZN => n229);
   U71 : INV_X1 port map( A => n32, ZN => n225);
   U72 : INV_X1 port map( A => n96, ZN => n194);
   U73 : INV_X1 port map( A => n34, ZN => n190);
   U74 : INV_X1 port map( A => n98, ZN => n230);
   U75 : INV_X1 port map( A => n36, ZN => n226);
   U76 : INV_X1 port map( A => n100, ZN => n195);
   U77 : INV_X1 port map( A => n38, ZN => n191);
   U78 : INV_X1 port map( A => n102, ZN => n231);
   U79 : INV_X1 port map( A => n40, ZN => n227);
   U80 : INV_X1 port map( A => n104, ZN => n183);
   U81 : INV_X1 port map( A => n42, ZN => n179);
   U82 : INV_X1 port map( A => n106, ZN => n219);
   U83 : INV_X1 port map( A => n44, ZN => n215);
   U84 : INV_X1 port map( A => n108, ZN => n184);
   U85 : INV_X1 port map( A => n46, ZN => n180);
   U86 : INV_X1 port map( A => n110, ZN => n220);
   U87 : INV_X1 port map( A => n48, ZN => n216);
   U88 : INV_X1 port map( A => n112, ZN => n185);
   U89 : INV_X1 port map( A => n50, ZN => n181);
   U90 : INV_X1 port map( A => n114, ZN => n221);
   U91 : INV_X1 port map( A => n52, ZN => n217);
   U92 : INV_X1 port map( A => n116, ZN => n186);
   U93 : INV_X1 port map( A => n54, ZN => n182);
   U94 : INV_X1 port map( A => n118, ZN => n222);
   U95 : INV_X1 port map( A => n56, ZN => n218);
   U96 : INV_X1 port map( A => n120, ZN => n201);
   U97 : INV_X1 port map( A => n58, ZN => n197);
   U98 : INV_X1 port map( A => n122, ZN => n237);
   U99 : INV_X1 port map( A => n60, ZN => n233);
   U100 : INV_X1 port map( A => n124, ZN => n202);
   U101 : INV_X1 port map( A => n62, ZN => n198);
   U102 : INV_X1 port map( A => n126, ZN => n238);
   U103 : INV_X1 port map( A => n64, ZN => n234);
   U104 : INV_X1 port map( A => n128, ZN => n203);
   U105 : INV_X1 port map( A => n66, ZN => n199);
   U106 : INV_X1 port map( A => n130, ZN => n239);
   U107 : INV_X1 port map( A => n68, ZN => n235);
   U108 : INV_X1 port map( A => n132, ZN => n204);
   U109 : INV_X1 port map( A => n70, ZN => n200);
   U110 : INV_X1 port map( A => n134, ZN => n240);
   U111 : INV_X1 port map( A => n72, ZN => n236);
   U112 : INV_X1 port map( A => n136, ZN => n177);
   U113 : INV_X1 port map( A => COARSE_38_port, ZN => n176);
   U114 : MUX2_X1 port map( A => COARSE_0_port, B => COARSE_4_port, S => 
                           DATA2(2), Z => n1);
   U115 : MUX2_X1 port map( A => n1, B => n170, S => DATA2(1), Z => n2);
   U116 : MUX2_X1 port map( A => n2, B => n206, S => DATA2(0), Z => 
                           SR_OUT_0_port);
   U117 : MUX2_X1 port map( A => n206, B => n169, S => DATA2(0), Z => 
                           SR_OUT_1_port);
   U118 : MUX2_X1 port map( A => n169, B => n207, S => DATA2(0), Z => 
                           SR_OUT_2_port);
   U119 : MUX2_X1 port map( A => n207, B => n171, S => DATA2(0), Z => 
                           SR_OUT_3_port);
   U120 : MUX2_X1 port map( A => n171, B => n208, S => DATA2(0), Z => 
                           SR_OUT_4_port);
   U121 : MUX2_X1 port map( A => n208, B => n172, S => DATA2(0), Z => 
                           SR_OUT_5_port);
   U122 : MUX2_X1 port map( A => n172, B => n209, S => DATA2(0), Z => 
                           SR_OUT_6_port);
   U123 : MUX2_X1 port map( A => n209, B => n188, S => DATA2(0), Z => 
                           SR_OUT_7_port);
   U124 : MUX2_X1 port map( A => n188, B => n224, S => DATA2(0), Z => 
                           SR_OUT_8_port);
   U125 : MUX2_X1 port map( A => n224, B => n189, S => DATA2(0), Z => 
                           SR_OUT_9_port);
   U126 : MUX2_X1 port map( A => n189, B => n225, S => DATA2(0), Z => 
                           SR_OUT_10_port);
   U127 : MUX2_X1 port map( A => n225, B => n190, S => DATA2(0), Z => 
                           SR_OUT_11_port);
   U128 : MUX2_X1 port map( A => n190, B => n226, S => DATA2(0), Z => 
                           SR_OUT_12_port);
   U129 : MUX2_X1 port map( A => n226, B => n191, S => DATA2(0), Z => 
                           SR_OUT_13_port);
   U130 : MUX2_X1 port map( A => n191, B => n227, S => DATA2(0), Z => 
                           SR_OUT_14_port);
   U131 : MUX2_X1 port map( A => n227, B => n179, S => DATA2(0), Z => 
                           SR_OUT_15_port);
   U132 : MUX2_X1 port map( A => n179, B => n215, S => DATA2(0), Z => 
                           SR_OUT_16_port);
   U133 : MUX2_X1 port map( A => n215, B => n180, S => DATA2(0), Z => 
                           SR_OUT_17_port);
   U134 : MUX2_X1 port map( A => n180, B => n216, S => DATA2(0), Z => 
                           SR_OUT_18_port);
   U135 : MUX2_X1 port map( A => n216, B => n181, S => DATA2(0), Z => 
                           SR_OUT_19_port);
   U136 : MUX2_X1 port map( A => n181, B => n217, S => DATA2(0), Z => 
                           SR_OUT_20_port);
   U137 : MUX2_X1 port map( A => n217, B => n182, S => DATA2(0), Z => 
                           SR_OUT_21_port);
   U138 : MUX2_X1 port map( A => n182, B => n218, S => DATA2(0), Z => 
                           SR_OUT_22_port);
   U139 : MUX2_X1 port map( A => n218, B => n197, S => DATA2(0), Z => 
                           SR_OUT_23_port);
   U140 : MUX2_X1 port map( A => n197, B => n233, S => DATA2(0), Z => 
                           SR_OUT_24_port);
   U141 : MUX2_X1 port map( A => n233, B => n198, S => DATA2(0), Z => 
                           SR_OUT_25_port);
   U142 : MUX2_X1 port map( A => n198, B => n234, S => DATA2(0), Z => 
                           SR_OUT_26_port);
   U143 : MUX2_X1 port map( A => n234, B => n199, S => DATA2(0), Z => 
                           SR_OUT_27_port);
   U144 : MUX2_X1 port map( A => n199, B => n235, S => DATA2(0), Z => 
                           SR_OUT_28_port);
   U145 : MUX2_X1 port map( A => n235, B => n200, S => DATA2(0), Z => 
                           SR_OUT_29_port);
   U146 : MUX2_X1 port map( A => n200, B => n236, S => DATA2(0), Z => 
                           SR_OUT_30_port);
   U147 : MUX2_X1 port map( A => COARSE_34_port, B => COARSE_38_port, S => 
                           DATA2(2), Z => n3);
   U148 : MUX2_X1 port map( A => n158, B => n3, S => DATA2(1), Z => n4);
   U149 : MUX2_X1 port map( A => n236, B => n4, S => DATA2(0), Z => 
                           SR_OUT_31_port);
   U150 : MUX2_X1 port map( A => COARSE_5_port, B => COARSE_1_port, S => 
                           DATA2(2), Z => n5);
   U151 : MUX2_X1 port map( A => n211, B => n5, S => DATA2(1), Z => n6);
   U152 : MUX2_X1 port map( A => n173, B => n6, S => DATA2(0), Z => 
                           SL_OUT_0_port);
   U153 : MUX2_X1 port map( A => n210, B => n173, S => DATA2(0), Z => 
                           SL_OUT_1_port);
   U154 : MUX2_X1 port map( A => n174, B => n210, S => DATA2(0), Z => 
                           SL_OUT_2_port);
   U155 : MUX2_X1 port map( A => n212, B => n174, S => DATA2(0), Z => 
                           SL_OUT_3_port);
   U156 : MUX2_X1 port map( A => n175, B => n212, S => DATA2(0), Z => 
                           SL_OUT_4_port);
   U157 : MUX2_X1 port map( A => n213, B => n175, S => DATA2(0), Z => 
                           SL_OUT_5_port);
   U158 : MUX2_X1 port map( A => n192, B => n213, S => DATA2(0), Z => 
                           SL_OUT_6_port);
   U159 : MUX2_X1 port map( A => n228, B => n192, S => DATA2(0), Z => 
                           SL_OUT_7_port);
   U160 : MUX2_X1 port map( A => n193, B => n228, S => DATA2(0), Z => 
                           SL_OUT_8_port);
   U161 : MUX2_X1 port map( A => n229, B => n193, S => DATA2(0), Z => 
                           SL_OUT_9_port);
   U162 : MUX2_X1 port map( A => n194, B => n229, S => DATA2(0), Z => 
                           SL_OUT_10_port);
   U163 : MUX2_X1 port map( A => n230, B => n194, S => DATA2(0), Z => 
                           SL_OUT_11_port);
   U164 : MUX2_X1 port map( A => n195, B => n230, S => DATA2(0), Z => 
                           SL_OUT_12_port);
   U165 : MUX2_X1 port map( A => n231, B => n195, S => DATA2(0), Z => 
                           SL_OUT_13_port);
   U166 : MUX2_X1 port map( A => n183, B => n231, S => DATA2(0), Z => 
                           SL_OUT_14_port);
   U167 : MUX2_X1 port map( A => n219, B => n183, S => DATA2(0), Z => 
                           SL_OUT_15_port);
   U168 : MUX2_X1 port map( A => n184, B => n219, S => DATA2(0), Z => 
                           SL_OUT_16_port);
   U169 : MUX2_X1 port map( A => n220, B => n184, S => DATA2(0), Z => 
                           SL_OUT_17_port);
   U170 : MUX2_X1 port map( A => n185, B => n220, S => DATA2(0), Z => 
                           SL_OUT_18_port);
   U171 : MUX2_X1 port map( A => n221, B => n185, S => DATA2(0), Z => 
                           SL_OUT_19_port);
   U172 : MUX2_X1 port map( A => n186, B => n221, S => DATA2(0), Z => 
                           SL_OUT_20_port);
   U173 : MUX2_X1 port map( A => n222, B => n186, S => DATA2(0), Z => 
                           SL_OUT_21_port);
   U174 : MUX2_X1 port map( A => n201, B => n222, S => DATA2(0), Z => 
                           SL_OUT_22_port);
   U175 : MUX2_X1 port map( A => n237, B => n201, S => DATA2(0), Z => 
                           SL_OUT_23_port);
   U176 : MUX2_X1 port map( A => n202, B => n237, S => DATA2(0), Z => 
                           SL_OUT_24_port);
   U177 : MUX2_X1 port map( A => n238, B => n202, S => DATA2(0), Z => 
                           SL_OUT_25_port);
   U178 : MUX2_X1 port map( A => n203, B => n238, S => DATA2(0), Z => 
                           SL_OUT_26_port);
   U179 : MUX2_X1 port map( A => n239, B => n203, S => DATA2(0), Z => 
                           SL_OUT_27_port);
   U180 : MUX2_X1 port map( A => n204, B => n239, S => DATA2(0), Z => 
                           SL_OUT_28_port);
   U181 : MUX2_X1 port map( A => n240, B => n204, S => DATA2(0), Z => 
                           SL_OUT_29_port);
   U182 : MUX2_X1 port map( A => n177, B => n240, S => DATA2(0), Z => 
                           SL_OUT_30_port);
   U183 : MUX2_X1 port map( A => COARSE_39_port, B => COARSE_35_port, S => 
                           DATA2(2), Z => n7);
   U184 : MUX2_X1 port map( A => n7, B => n164, S => DATA2(1), Z => n8);
   U185 : MUX2_X1 port map( A => n8, B => n177, S => DATA2(0), Z => 
                           SL_OUT_31_port);
   U186 : MUX2_X1 port map( A => n151, B => n205, S => DATA2(2), Z => n9);
   U187 : MUX2_X1 port map( A => n143, B => n162, S => DATA2(2), Z => n10);
   U188 : MUX2_X1 port map( A => n10, B => n9, S => DATA2(1), Z => n11);
   U189 : MUX2_X1 port map( A => n147, B => n168, S => DATA2(2), Z => n12);
   U190 : MUX2_X1 port map( A => n156, B => n137, S => DATA2(2), Z => n13);
   U191 : MUX2_X1 port map( A => n12, B => n13, S => DATA2(1), Z => n14);
   U192 : MUX2_X1 port map( A => n162, B => n141, S => DATA2(2), Z => n15);
   U193 : MUX2_X1 port map( A => n9, B => n15, S => DATA2(1), Z => n16);
   U194 : MUX2_X1 port map( A => n168, B => n149, S => DATA2(2), Z => n17);
   U195 : MUX2_X1 port map( A => n13, B => n17, S => DATA2(1), Z => n18);
   U196 : MUX2_X1 port map( A => n205, B => n154, S => DATA2(2), Z => n19);
   U197 : MUX2_X1 port map( A => n15, B => n19, S => DATA2(1), Z => n20);
   U198 : MUX2_X1 port map( A => n137, B => n160, S => DATA2(2), Z => n21);
   U199 : MUX2_X1 port map( A => n17, B => n21, S => DATA2(1), Z => n22);
   U200 : MUX2_X1 port map( A => n141, B => n166, S => DATA2(2), Z => n23);
   U201 : MUX2_X1 port map( A => n19, B => n23, S => DATA2(1), Z => n24);
   U202 : MUX2_X1 port map( A => n149, B => n187, S => DATA2(2), Z => n25);
   U203 : MUX2_X1 port map( A => n21, B => n25, S => DATA2(1), Z => n26);
   U204 : MUX2_X1 port map( A => n154, B => n223, S => DATA2(2), Z => n27);
   U205 : MUX2_X1 port map( A => n23, B => n27, S => DATA2(1), Z => n28);
   U206 : MUX2_X1 port map( A => n160, B => n139, S => DATA2(2), Z => n29);
   U207 : MUX2_X1 port map( A => n25, B => n29, S => DATA2(1), Z => n30);
   U208 : MUX2_X1 port map( A => n166, B => n144, S => DATA2(2), Z => n31);
   U209 : MUX2_X1 port map( A => n27, B => n31, S => DATA2(1), Z => n32);
   U210 : MUX2_X1 port map( A => n187, B => n148, S => DATA2(2), Z => n33);
   U211 : MUX2_X1 port map( A => n29, B => n33, S => DATA2(1), Z => n34);
   U212 : MUX2_X1 port map( A => n223, B => n153, S => DATA2(2), Z => n35);
   U213 : MUX2_X1 port map( A => n31, B => n35, S => DATA2(1), Z => n36);
   U214 : MUX2_X1 port map( A => n139, B => n159, S => DATA2(2), Z => n37);
   U215 : MUX2_X1 port map( A => n33, B => n37, S => DATA2(1), Z => n38);
   U216 : MUX2_X1 port map( A => n144, B => n165, S => DATA2(2), Z => n39);
   U217 : MUX2_X1 port map( A => n35, B => n39, S => DATA2(1), Z => n40);
   U218 : MUX2_X1 port map( A => n148, B => n178, S => DATA2(2), Z => n41);
   U219 : MUX2_X1 port map( A => n37, B => n41, S => DATA2(1), Z => n42);
   U220 : MUX2_X1 port map( A => n153, B => n214, S => DATA2(2), Z => n43);
   U221 : MUX2_X1 port map( A => n39, B => n43, S => DATA2(1), Z => n44);
   U222 : MUX2_X1 port map( A => n159, B => n140, S => DATA2(2), Z => n45);
   U223 : MUX2_X1 port map( A => n41, B => n45, S => DATA2(1), Z => n46);
   U224 : MUX2_X1 port map( A => n165, B => n145, S => DATA2(2), Z => n47);
   U225 : MUX2_X1 port map( A => n43, B => n47, S => DATA2(1), Z => n48);
   U226 : MUX2_X1 port map( A => n178, B => n150, S => DATA2(2), Z => n49);
   U227 : MUX2_X1 port map( A => n45, B => n49, S => DATA2(1), Z => n50);
   U228 : MUX2_X1 port map( A => n214, B => n155, S => DATA2(2), Z => n51);
   U229 : MUX2_X1 port map( A => n47, B => n51, S => DATA2(1), Z => n52);
   U230 : MUX2_X1 port map( A => n140, B => n161, S => DATA2(2), Z => n53);
   U231 : MUX2_X1 port map( A => n49, B => n53, S => DATA2(1), Z => n54);
   U232 : MUX2_X1 port map( A => n145, B => n167, S => DATA2(2), Z => n55);
   U233 : MUX2_X1 port map( A => n51, B => n55, S => DATA2(1), Z => n56);
   U234 : MUX2_X1 port map( A => n150, B => n196, S => DATA2(2), Z => n57);
   U235 : MUX2_X1 port map( A => n53, B => n57, S => DATA2(1), Z => n58);
   U236 : MUX2_X1 port map( A => n155, B => n232, S => DATA2(2), Z => n59);
   U237 : MUX2_X1 port map( A => n55, B => n59, S => DATA2(1), Z => n60);
   U238 : MUX2_X1 port map( A => n161, B => n138, S => DATA2(2), Z => n61);
   U239 : MUX2_X1 port map( A => n57, B => n61, S => DATA2(1), Z => n62);
   U240 : MUX2_X1 port map( A => n167, B => n142, S => DATA2(2), Z => n63);
   U241 : MUX2_X1 port map( A => n59, B => n63, S => DATA2(1), Z => n64);
   U242 : MUX2_X1 port map( A => n196, B => n146, S => DATA2(2), Z => n65);
   U243 : MUX2_X1 port map( A => n61, B => n65, S => DATA2(1), Z => n66);
   U244 : MUX2_X1 port map( A => n232, B => n152, S => DATA2(2), Z => n67);
   U245 : MUX2_X1 port map( A => n63, B => n67, S => DATA2(1), Z => n68);
   U246 : MUX2_X1 port map( A => n138, B => n157, S => DATA2(2), Z => n69);
   U247 : MUX2_X1 port map( A => n65, B => n69, S => DATA2(1), Z => n70);
   U248 : MUX2_X1 port map( A => n142, B => n163, S => DATA2(2), Z => n71);
   U249 : MUX2_X1 port map( A => n67, B => n71, S => DATA2(1), Z => n72);
   U250 : MUX2_X1 port map( A => n205, B => n151, S => DATA2(2), Z => n73);
   U251 : MUX2_X1 port map( A => n168, B => n147, S => DATA2(2), Z => n74);
   U252 : MUX2_X1 port map( A => n137, B => n156, S => DATA2(2), Z => n75);
   U253 : MUX2_X1 port map( A => n75, B => n74, S => DATA2(1), Z => n76);
   U254 : MUX2_X1 port map( A => n141, B => n162, S => DATA2(2), Z => n77);
   U255 : MUX2_X1 port map( A => n77, B => n73, S => DATA2(1), Z => n78);
   U256 : MUX2_X1 port map( A => n149, B => n168, S => DATA2(2), Z => n79);
   U257 : MUX2_X1 port map( A => n79, B => n75, S => DATA2(1), Z => n80);
   U258 : MUX2_X1 port map( A => n154, B => n205, S => DATA2(2), Z => n81);
   U259 : MUX2_X1 port map( A => n81, B => n77, S => DATA2(1), Z => n82);
   U260 : MUX2_X1 port map( A => n160, B => n137, S => DATA2(2), Z => n83);
   U261 : MUX2_X1 port map( A => n83, B => n79, S => DATA2(1), Z => n84);
   U262 : MUX2_X1 port map( A => n166, B => n141, S => DATA2(2), Z => n85);
   U263 : MUX2_X1 port map( A => n85, B => n81, S => DATA2(1), Z => n86);
   U264 : MUX2_X1 port map( A => n187, B => n149, S => DATA2(2), Z => n87);
   U265 : MUX2_X1 port map( A => n87, B => n83, S => DATA2(1), Z => n88);
   U266 : MUX2_X1 port map( A => n223, B => n154, S => DATA2(2), Z => n89);
   U267 : MUX2_X1 port map( A => n89, B => n85, S => DATA2(1), Z => n90);
   U268 : MUX2_X1 port map( A => n139, B => n160, S => DATA2(2), Z => n91);
   U269 : MUX2_X1 port map( A => n91, B => n87, S => DATA2(1), Z => n92);
   U270 : MUX2_X1 port map( A => n144, B => n166, S => DATA2(2), Z => n93);
   U271 : MUX2_X1 port map( A => n93, B => n89, S => DATA2(1), Z => n94);
   U272 : MUX2_X1 port map( A => n148, B => n187, S => DATA2(2), Z => n95);
   U273 : MUX2_X1 port map( A => n95, B => n91, S => DATA2(1), Z => n96);
   U274 : MUX2_X1 port map( A => n153, B => n223, S => DATA2(2), Z => n97);
   U275 : MUX2_X1 port map( A => n97, B => n93, S => DATA2(1), Z => n98);
   U276 : MUX2_X1 port map( A => n159, B => n139, S => DATA2(2), Z => n99);
   U277 : MUX2_X1 port map( A => n99, B => n95, S => DATA2(1), Z => n100);
   U278 : MUX2_X1 port map( A => n165, B => n144, S => DATA2(2), Z => n101);
   U279 : MUX2_X1 port map( A => n101, B => n97, S => DATA2(1), Z => n102);
   U280 : MUX2_X1 port map( A => n178, B => n148, S => DATA2(2), Z => n103);
   U281 : MUX2_X1 port map( A => n103, B => n99, S => DATA2(1), Z => n104);
   U282 : MUX2_X1 port map( A => n214, B => n153, S => DATA2(2), Z => n105);
   U283 : MUX2_X1 port map( A => n105, B => n101, S => DATA2(1), Z => n106);
   U284 : MUX2_X1 port map( A => n140, B => n159, S => DATA2(2), Z => n107);
   U285 : MUX2_X1 port map( A => n107, B => n103, S => DATA2(1), Z => n108);
   U286 : MUX2_X1 port map( A => n145, B => n165, S => DATA2(2), Z => n109);
   U287 : MUX2_X1 port map( A => n109, B => n105, S => DATA2(1), Z => n110);
   U288 : MUX2_X1 port map( A => n150, B => n178, S => DATA2(2), Z => n111);
   U289 : MUX2_X1 port map( A => n111, B => n107, S => DATA2(1), Z => n112);
   U290 : MUX2_X1 port map( A => n155, B => n214, S => DATA2(2), Z => n113);
   U291 : MUX2_X1 port map( A => n113, B => n109, S => DATA2(1), Z => n114);
   U292 : MUX2_X1 port map( A => n161, B => n140, S => DATA2(2), Z => n115);
   U293 : MUX2_X1 port map( A => n115, B => n111, S => DATA2(1), Z => n116);
   U294 : MUX2_X1 port map( A => n167, B => n145, S => DATA2(2), Z => n117);
   U295 : MUX2_X1 port map( A => n117, B => n113, S => DATA2(1), Z => n118);
   U296 : MUX2_X1 port map( A => n196, B => n150, S => DATA2(2), Z => n119);
   U297 : MUX2_X1 port map( A => n119, B => n115, S => DATA2(1), Z => n120);
   U298 : MUX2_X1 port map( A => n232, B => n155, S => DATA2(2), Z => n121);
   U299 : MUX2_X1 port map( A => n121, B => n117, S => DATA2(1), Z => n122);
   U300 : MUX2_X1 port map( A => n138, B => n161, S => DATA2(2), Z => n123);
   U301 : MUX2_X1 port map( A => n123, B => n119, S => DATA2(1), Z => n124);
   U302 : MUX2_X1 port map( A => n142, B => n167, S => DATA2(2), Z => n125);
   U303 : MUX2_X1 port map( A => n125, B => n121, S => DATA2(1), Z => n126);
   U304 : MUX2_X1 port map( A => n146, B => n196, S => DATA2(2), Z => n127);
   U305 : MUX2_X1 port map( A => n127, B => n123, S => DATA2(1), Z => n128);
   U306 : MUX2_X1 port map( A => n152, B => n232, S => DATA2(2), Z => n129);
   U307 : MUX2_X1 port map( A => n129, B => n125, S => DATA2(1), Z => n130);
   U308 : MUX2_X1 port map( A => n157, B => n138, S => DATA2(2), Z => n131);
   U309 : MUX2_X1 port map( A => n131, B => n127, S => DATA2(1), Z => n132);
   U310 : MUX2_X1 port map( A => n163, B => n142, S => DATA2(2), Z => n133);
   U311 : MUX2_X1 port map( A => n133, B => n129, S => DATA2(1), Z => n134);
   U312 : MUX2_X1 port map( A => n176, B => n146, S => DATA2(2), Z => n135);
   U313 : MUX2_X1 port map( A => n135, B => n131, S => DATA2(1), Z => n136);
   U314 : MUX2_X1 port map( A => SR_OUT_30_port, B => SL_OUT_30_port, S => n241
                           , Z => OUTPUT(30));
   U315 : MUX2_X1 port map( A => SR_OUT_29_port, B => SL_OUT_29_port, S => n241
                           , Z => OUTPUT(29));
   U316 : MUX2_X1 port map( A => SR_OUT_28_port, B => SL_OUT_28_port, S => n241
                           , Z => OUTPUT(28));
   U317 : MUX2_X1 port map( A => SR_OUT_27_port, B => SL_OUT_27_port, S => n241
                           , Z => OUTPUT(27));
   U318 : MUX2_X1 port map( A => SR_OUT_26_port, B => SL_OUT_26_port, S => n241
                           , Z => OUTPUT(26));
   U319 : MUX2_X1 port map( A => SR_OUT_25_port, B => SL_OUT_25_port, S => n241
                           , Z => OUTPUT(25));
   U320 : MUX2_X1 port map( A => SR_OUT_24_port, B => SL_OUT_24_port, S => n241
                           , Z => OUTPUT(24));
   U321 : MUX2_X1 port map( A => SR_OUT_23_port, B => SL_OUT_23_port, S => n241
                           , Z => OUTPUT(23));
   U322 : MUX2_X1 port map( A => SR_OUT_31_port, B => SL_OUT_31_port, S => n241
                           , Z => OUTPUT(31));
   U323 : MUX2_X1 port map( A => SR_OUT_14_port, B => SL_OUT_14_port, S => n241
                           , Z => OUTPUT(14));
   U324 : MUX2_X1 port map( A => SR_OUT_13_port, B => SL_OUT_13_port, S => n241
                           , Z => OUTPUT(13));
   U325 : MUX2_X1 port map( A => SR_OUT_12_port, B => SL_OUT_12_port, S => n241
                           , Z => OUTPUT(12));
   U326 : MUX2_X1 port map( A => SR_OUT_11_port, B => SL_OUT_11_port, S => n241
                           , Z => OUTPUT(11));
   U327 : MUX2_X1 port map( A => SR_OUT_10_port, B => SL_OUT_10_port, S => n241
                           , Z => OUTPUT(10));
   U328 : MUX2_X1 port map( A => SR_OUT_9_port, B => SL_OUT_9_port, S => n241, 
                           Z => OUTPUT(9));
   U329 : MUX2_X1 port map( A => SR_OUT_8_port, B => SL_OUT_8_port, S => n241, 
                           Z => OUTPUT(8));
   U330 : MUX2_X1 port map( A => SR_OUT_7_port, B => SL_OUT_7_port, S => n241, 
                           Z => OUTPUT(7));
   U331 : MUX2_X1 port map( A => SR_OUT_15_port, B => SL_OUT_15_port, S => n241
                           , Z => OUTPUT(15));
   U332 : MUX2_X1 port map( A => SR_OUT_22_port, B => SL_OUT_22_port, S => n241
                           , Z => OUTPUT(22));
   U333 : MUX2_X1 port map( A => SR_OUT_21_port, B => SL_OUT_21_port, S => n241
                           , Z => OUTPUT(21));
   U334 : MUX2_X1 port map( A => SR_OUT_20_port, B => SL_OUT_20_port, S => n241
                           , Z => OUTPUT(20));
   U335 : MUX2_X1 port map( A => SR_OUT_19_port, B => SL_OUT_19_port, S => n241
                           , Z => OUTPUT(19));
   U336 : MUX2_X1 port map( A => SR_OUT_18_port, B => SL_OUT_18_port, S => n241
                           , Z => OUTPUT(18));
   U337 : MUX2_X1 port map( A => SR_OUT_17_port, B => SL_OUT_17_port, S => n241
                           , Z => OUTPUT(17));
   U338 : MUX2_X1 port map( A => SR_OUT_16_port, B => SL_OUT_16_port, S => n241
                           , Z => OUTPUT(16));
   U339 : MUX2_X1 port map( A => SR_OUT_6_port, B => SL_OUT_6_port, S => n241, 
                           Z => OUTPUT(6));
   U340 : MUX2_X1 port map( A => SR_OUT_5_port, B => SL_OUT_5_port, S => n241, 
                           Z => OUTPUT(5));
   U341 : MUX2_X1 port map( A => SR_OUT_4_port, B => SL_OUT_4_port, S => n241, 
                           Z => OUTPUT(4));
   U342 : MUX2_X1 port map( A => SR_OUT_3_port, B => SL_OUT_3_port, S => n241, 
                           Z => OUTPUT(3));
   U343 : MUX2_X1 port map( A => SR_OUT_0_port, B => SL_OUT_0_port, S => n241, 
                           Z => OUTPUT(0));
   U344 : MUX2_X1 port map( A => SR_OUT_2_port, B => SL_OUT_2_port, S => n241, 
                           Z => OUTPUT(2));
   U345 : MUX2_X1 port map( A => SR_OUT_1_port, B => SL_OUT_1_port, S => n241, 
                           Z => OUTPUT(1));
   U346 : OAI221_X1 port map( B1 => n242, B2 => n243, C1 => n244, C2 => n245, A
                           => n246, ZN => COARSE_9_port);
   U347 : AOI22_X1 port map( A1 => DATA1(1), A2 => n247, B1 => DATA1(25), B2 =>
                           n248, ZN => n246);
   U348 : OAI221_X1 port map( B1 => n242, B2 => n249, C1 => n244, C2 => n250, A
                           => n251, ZN => COARSE_8_port);
   U349 : AOI22_X1 port map( A1 => DATA1(0), A2 => n247, B1 => DATA1(24), B2 =>
                           n248, ZN => n251);
   U350 : OAI221_X1 port map( B1 => n242, B2 => n252, C1 => n244, C2 => n253, A
                           => n254, ZN => COARSE_7_port);
   U351 : AOI22_X1 port map( A1 => DATA1(23), A2 => n248, B1 => DATA1(31), B2 
                           => n255, ZN => n254);
   U352 : INV_X1 port map( A => DATA1(7), ZN => n252);
   U353 : OAI221_X1 port map( B1 => n242, B2 => n256, C1 => n244, C2 => n257, A
                           => n258, ZN => COARSE_6_port);
   U354 : AOI22_X1 port map( A1 => DATA1(22), A2 => n248, B1 => DATA1(30), B2 
                           => n255, ZN => n258);
   U355 : INV_X1 port map( A => DATA1(6), ZN => n256);
   U356 : OAI221_X1 port map( B1 => n242, B2 => n259, C1 => n244, C2 => n260, A
                           => n261, ZN => COARSE_5_port);
   U357 : AOI22_X1 port map( A1 => DATA1(21), A2 => n248, B1 => DATA1(29), B2 
                           => n255, ZN => n261);
   U358 : INV_X1 port map( A => DATA1(5), ZN => n259);
   U359 : OAI221_X1 port map( B1 => n242, B2 => n262, C1 => n244, C2 => n263, A
                           => n264, ZN => COARSE_4_port);
   U360 : AOI22_X1 port map( A1 => DATA1(20), A2 => n248, B1 => DATA1(28), B2 
                           => n255, ZN => n264);
   U361 : INV_X1 port map( A => DATA1(4), ZN => n262);
   U362 : OAI221_X1 port map( B1 => n242, B2 => n265, C1 => n244, C2 => n266, A
                           => n267, ZN => COARSE_3_port);
   U363 : AOI22_X1 port map( A1 => DATA1(19), A2 => n248, B1 => DATA1(27), B2 
                           => n255, ZN => n267);
   U364 : INV_X1 port map( A => DATA1(3), ZN => n265);
   U365 : OAI221_X1 port map( B1 => n268, B2 => n269, C1 => n270, C2 => n271, A
                           => n272, ZN => COARSE_39_port);
   U366 : AOI22_X1 port map( A1 => n273, A2 => DATA1(7), B1 => n274, B2 => 
                           DATA1(15), ZN => n272);
   U367 : OAI221_X1 port map( B1 => n275, B2 => n269, C1 => n270, C2 => n276, A
                           => n277, ZN => COARSE_38_port);
   U368 : AOI22_X1 port map( A1 => n273, A2 => DATA1(6), B1 => n274, B2 => 
                           DATA1(14), ZN => n277);
   U369 : OAI221_X1 port map( B1 => n278, B2 => n269, C1 => n270, C2 => n279, A
                           => n280, ZN => COARSE_37_port);
   U370 : AOI22_X1 port map( A1 => n273, A2 => DATA1(5), B1 => n274, B2 => 
                           DATA1(13), ZN => n280);
   U371 : OAI221_X1 port map( B1 => n281, B2 => n269, C1 => n270, C2 => n282, A
                           => n283, ZN => COARSE_36_port);
   U372 : AOI22_X1 port map( A1 => n273, A2 => DATA1(4), B1 => n274, B2 => 
                           DATA1(12), ZN => n283);
   U373 : OAI221_X1 port map( B1 => n284, B2 => n269, C1 => n270, C2 => n285, A
                           => n286, ZN => COARSE_35_port);
   U374 : AOI22_X1 port map( A1 => n273, A2 => DATA1(3), B1 => n274, B2 => 
                           DATA1(11), ZN => n286);
   U375 : OAI221_X1 port map( B1 => n269, B2 => n287, C1 => n270, C2 => n288, A
                           => n289, ZN => COARSE_34_port);
   U376 : AOI22_X1 port map( A1 => DATA1(2), A2 => n273, B1 => DATA1(10), B2 =>
                           n274, ZN => n289);
   U377 : OAI221_X1 port map( B1 => n245, B2 => n269, C1 => n270, C2 => n290, A
                           => n291, ZN => COARSE_33_port);
   U378 : AOI22_X1 port map( A1 => n273, A2 => DATA1(1), B1 => n274, B2 => 
                           DATA1(9), ZN => n291);
   U379 : OAI221_X1 port map( B1 => n250, B2 => n269, C1 => n270, C2 => n292, A
                           => n293, ZN => COARSE_32_port);
   U380 : AOI22_X1 port map( A1 => n273, A2 => DATA1(0), B1 => n274, B2 => 
                           DATA1(8), ZN => n293);
   U381 : INV_X1 port map( A => n296, ZN => n269);
   U382 : OAI221_X1 port map( B1 => n270, B2 => n268, C1 => n242, C2 => n271, A
                           => n297, ZN => COARSE_31_port);
   U383 : AOI22_X1 port map( A1 => n274, A2 => DATA1(7), B1 => n296, B2 => 
                           DATA1(15), ZN => n297);
   U384 : OAI221_X1 port map( B1 => n270, B2 => n275, C1 => n242, C2 => n276, A
                           => n298, ZN => COARSE_30_port);
   U385 : AOI22_X1 port map( A1 => n274, A2 => DATA1(6), B1 => n296, B2 => 
                           DATA1(14), ZN => n298);
   U386 : OAI221_X1 port map( B1 => n242, B2 => n299, C1 => n244, C2 => n300, A
                           => n301, ZN => COARSE_2_port);
   U387 : AOI22_X1 port map( A1 => DATA1(18), A2 => n248, B1 => DATA1(26), B2 
                           => n255, ZN => n301);
   U388 : INV_X1 port map( A => DATA1(2), ZN => n299);
   U389 : OAI221_X1 port map( B1 => n270, B2 => n278, C1 => n242, C2 => n279, A
                           => n302, ZN => COARSE_29_port);
   U390 : AOI22_X1 port map( A1 => n274, A2 => DATA1(5), B1 => n296, B2 => 
                           DATA1(13), ZN => n302);
   U391 : OAI221_X1 port map( B1 => n270, B2 => n281, C1 => n242, C2 => n282, A
                           => n303, ZN => COARSE_28_port);
   U392 : AOI22_X1 port map( A1 => n274, A2 => DATA1(4), B1 => n296, B2 => 
                           DATA1(12), ZN => n303);
   U393 : OAI221_X1 port map( B1 => n270, B2 => n284, C1 => n242, C2 => n285, A
                           => n304, ZN => COARSE_27_port);
   U394 : AOI22_X1 port map( A1 => n274, A2 => DATA1(3), B1 => n296, B2 => 
                           DATA1(11), ZN => n304);
   U395 : OAI221_X1 port map( B1 => n270, B2 => n287, C1 => n242, C2 => n288, A
                           => n305, ZN => COARSE_26_port);
   U396 : AOI22_X1 port map( A1 => DATA1(2), A2 => n274, B1 => DATA1(10), B2 =>
                           n296, ZN => n305);
   U397 : OAI221_X1 port map( B1 => n270, B2 => n245, C1 => n290, C2 => n242, A
                           => n306, ZN => COARSE_25_port);
   U398 : AOI22_X1 port map( A1 => n274, A2 => DATA1(1), B1 => n296, B2 => 
                           DATA1(9), ZN => n306);
   U399 : OAI221_X1 port map( B1 => n270, B2 => n250, C1 => n242, C2 => n292, A
                           => n307, ZN => COARSE_24_port);
   U400 : AOI22_X1 port map( A1 => n274, A2 => DATA1(0), B1 => n296, B2 => 
                           DATA1(8), ZN => n307);
   U401 : INV_X1 port map( A => n247, ZN => n270);
   U402 : OAI221_X1 port map( B1 => n242, B2 => n268, C1 => n244, C2 => n271, A
                           => n308, ZN => COARSE_23_port);
   U403 : AOI22_X1 port map( A1 => n296, A2 => DATA1(7), B1 => DATA1(15), B2 =>
                           n247, ZN => n308);
   U404 : INV_X1 port map( A => DATA1(31), ZN => n271);
   U405 : OAI221_X1 port map( B1 => n242, B2 => n275, C1 => n244, C2 => n276, A
                           => n309, ZN => COARSE_22_port);
   U406 : AOI22_X1 port map( A1 => n296, A2 => DATA1(6), B1 => DATA1(14), B2 =>
                           n247, ZN => n309);
   U407 : INV_X1 port map( A => DATA1(30), ZN => n276);
   U408 : OAI221_X1 port map( B1 => n242, B2 => n278, C1 => n244, C2 => n279, A
                           => n310, ZN => COARSE_21_port);
   U409 : AOI22_X1 port map( A1 => n296, A2 => DATA1(5), B1 => DATA1(13), B2 =>
                           n247, ZN => n310);
   U410 : INV_X1 port map( A => DATA1(29), ZN => n279);
   U411 : OAI221_X1 port map( B1 => n242, B2 => n281, C1 => n244, C2 => n282, A
                           => n311, ZN => COARSE_20_port);
   U412 : AOI22_X1 port map( A1 => n296, A2 => DATA1(4), B1 => DATA1(12), B2 =>
                           n247, ZN => n311);
   U413 : INV_X1 port map( A => DATA1(28), ZN => n282);
   U414 : OAI221_X1 port map( B1 => n312, B2 => n242, C1 => n243, C2 => n244, A
                           => n313, ZN => COARSE_1_port);
   U415 : AOI22_X1 port map( A1 => DATA1(17), A2 => n248, B1 => n255, B2 => 
                           DATA1(25), ZN => n313);
   U416 : INV_X1 port map( A => DATA1(9), ZN => n243);
   U417 : INV_X1 port map( A => DATA1(1), ZN => n312);
   U418 : OAI221_X1 port map( B1 => n242, B2 => n284, C1 => n244, C2 => n285, A
                           => n314, ZN => COARSE_19_port);
   U419 : AOI22_X1 port map( A1 => n296, A2 => DATA1(3), B1 => DATA1(11), B2 =>
                           n247, ZN => n314);
   U420 : INV_X1 port map( A => DATA1(27), ZN => n285);
   U421 : OAI221_X1 port map( B1 => n242, B2 => n287, C1 => n244, C2 => n288, A
                           => n315, ZN => COARSE_18_port);
   U422 : AOI22_X1 port map( A1 => DATA1(2), A2 => n296, B1 => DATA1(10), B2 =>
                           n247, ZN => n315);
   U423 : INV_X1 port map( A => DATA1(26), ZN => n288);
   U424 : OAI221_X1 port map( B1 => n242, B2 => n245, C1 => n290, C2 => n244, A
                           => n316, ZN => COARSE_17_port);
   U425 : AOI22_X1 port map( A1 => n296, A2 => DATA1(1), B1 => DATA1(9), B2 => 
                           n247, ZN => n316);
   U426 : INV_X1 port map( A => DATA1(25), ZN => n290);
   U427 : INV_X1 port map( A => DATA1(17), ZN => n245);
   U428 : OAI221_X1 port map( B1 => n242, B2 => n250, C1 => n244, C2 => n292, A
                           => n317, ZN => COARSE_16_port);
   U429 : AOI22_X1 port map( A1 => n296, A2 => DATA1(0), B1 => DATA1(8), B2 => 
                           n247, ZN => n317);
   U430 : INV_X1 port map( A => DATA1(24), ZN => n292);
   U431 : INV_X1 port map( A => DATA1(16), ZN => n250);
   U432 : OAI221_X1 port map( B1 => n242, B2 => n253, C1 => n244, C2 => n268, A
                           => n318, ZN => COARSE_15_port);
   U433 : AOI22_X1 port map( A1 => DATA1(7), A2 => n247, B1 => DATA1(31), B2 =>
                           n248, ZN => n318);
   U434 : INV_X1 port map( A => DATA1(23), ZN => n268);
   U435 : INV_X1 port map( A => DATA1(15), ZN => n253);
   U436 : OAI221_X1 port map( B1 => n242, B2 => n257, C1 => n244, C2 => n275, A
                           => n319, ZN => COARSE_14_port);
   U437 : AOI22_X1 port map( A1 => DATA1(6), A2 => n247, B1 => DATA1(30), B2 =>
                           n248, ZN => n319);
   U438 : INV_X1 port map( A => DATA1(22), ZN => n275);
   U439 : INV_X1 port map( A => DATA1(14), ZN => n257);
   U440 : OAI221_X1 port map( B1 => n242, B2 => n260, C1 => n244, C2 => n278, A
                           => n320, ZN => COARSE_13_port);
   U441 : AOI22_X1 port map( A1 => DATA1(5), A2 => n247, B1 => DATA1(29), B2 =>
                           n248, ZN => n320);
   U442 : INV_X1 port map( A => DATA1(21), ZN => n278);
   U443 : INV_X1 port map( A => DATA1(13), ZN => n260);
   U444 : OAI221_X1 port map( B1 => n242, B2 => n263, C1 => n244, C2 => n281, A
                           => n321, ZN => COARSE_12_port);
   U445 : AOI22_X1 port map( A1 => DATA1(4), A2 => n247, B1 => DATA1(28), B2 =>
                           n248, ZN => n321);
   U446 : INV_X1 port map( A => DATA1(20), ZN => n281);
   U447 : INV_X1 port map( A => DATA1(12), ZN => n263);
   U448 : OAI221_X1 port map( B1 => n242, B2 => n266, C1 => n244, C2 => n284, A
                           => n322, ZN => COARSE_11_port);
   U449 : AOI22_X1 port map( A1 => DATA1(3), A2 => n247, B1 => DATA1(27), B2 =>
                           n248, ZN => n322);
   U450 : INV_X1 port map( A => DATA1(19), ZN => n284);
   U451 : INV_X1 port map( A => DATA1(11), ZN => n266);
   U452 : OAI221_X1 port map( B1 => n242, B2 => n300, C1 => n244, C2 => n287, A
                           => n323, ZN => COARSE_10_port);
   U453 : AOI22_X1 port map( A1 => DATA1(2), A2 => n247, B1 => DATA1(26), B2 =>
                           n248, ZN => n323);
   U454 : INV_X1 port map( A => DATA1(18), ZN => n287);
   U455 : INV_X1 port map( A => DATA1(10), ZN => n300);
   U456 : OAI221_X1 port map( B1 => n242, B2 => n324, C1 => n244, C2 => n249, A
                           => n325, ZN => COARSE_0_port);
   U457 : AOI22_X1 port map( A1 => DATA1(16), A2 => n248, B1 => n255, B2 => 
                           DATA1(24), ZN => n325);
   U458 : INV_X1 port map( A => DATA1(8), ZN => n249);
   U459 : NAND3_X1 port map( A1 => CONF, A2 => n294, A3 => DATA2(3), ZN => n244
                           );
   U460 : INV_X1 port map( A => DATA1(0), ZN => n324);
   U461 : INV_X1 port map( A => DATA2(4), ZN => n294);
   U462 : INV_X1 port map( A => DATA2(3), ZN => n295);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_0 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_0;

architecture SYN_BEHAVIOUR of NAND4_0 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_0 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_0;

architecture SYN_BEHAVIOUR of NAND3_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32 is

   port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
         downto 0));

end ALU_N32;

architecture SYN_BEHAVIOR of ALU_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ALU_N32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component ALU_N32_DW01_addsub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (31 downto 0);  CO : out 
            std_logic);
   end component;
   
   component BARREL_SHIFTER_N32
      port( CONF : in std_logic;  DATA1, DATA2 : in std_logic_vector (31 downto
            0);  OUTPUT : out std_logic_vector (31 downto 0));
   end component;
   
   component NAND4_1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_2
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_3
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_4
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_5
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_6
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_7
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_8
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_9
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_10
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_11
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_12
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_13
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_14
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_15
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_16
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_17
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_18
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_19
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_20
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_21
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_22
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_23
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_24
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_25
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_26
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_27
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_28
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_29
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_30
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_31
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_0
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_2
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_3
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_4
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_5
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_6
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_7
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_8
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_9
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_10
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_11
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_12
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_13
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_14
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_15
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_16
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_17
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_18
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_19
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_20
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_21
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_22
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_23
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_24
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_25
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_26
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_27
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_28
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_29
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_30
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_31
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_32
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_33
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_34
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_35
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_36
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_37
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_38
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_39
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_40
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_41
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_42
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_43
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_44
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_45
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_46
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_47
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_48
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_49
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_50
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_51
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_52
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_53
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_54
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_55
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_56
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_57
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_58
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_59
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_60
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_61
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_62
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_63
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_64
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_65
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_66
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_67
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_68
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_69
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_70
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_71
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_72
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_73
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_74
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_75
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_76
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_77
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_78
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_79
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_80
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_81
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_82
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_83
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_84
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_85
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_86
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_87
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_88
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_89
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_90
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_91
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_92
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_93
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_94
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_95
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_96
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_97
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_98
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_99
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_100
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_101
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_102
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_103
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_104
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_105
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_106
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_107
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_108
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_109
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_110
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_111
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_112
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_113
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_114
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_115
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_116
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_117
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_118
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_119
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_120
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_121
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_122
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_123
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_124
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_125
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_126
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_127
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_0
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89,
      N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
      N104, N105, N106, N107, N108, N109, N110, Y_LOGIC_31_port, 
      Y_LOGIC_30_port, Y_LOGIC_29_port, Y_LOGIC_28_port, Y_LOGIC_27_port, 
      Y_LOGIC_26_port, Y_LOGIC_25_port, Y_LOGIC_24_port, Y_LOGIC_23_port, 
      Y_LOGIC_22_port, Y_LOGIC_21_port, Y_LOGIC_20_port, Y_LOGIC_19_port, 
      Y_LOGIC_18_port, Y_LOGIC_17_port, Y_LOGIC_16_port, Y_LOGIC_15_port, 
      Y_LOGIC_14_port, Y_LOGIC_13_port, Y_LOGIC_12_port, Y_LOGIC_11_port, 
      Y_LOGIC_10_port, Y_LOGIC_9_port, Y_LOGIC_8_port, Y_LOGIC_7_port, 
      Y_LOGIC_6_port, Y_LOGIC_5_port, Y_LOGIC_4_port, Y_LOGIC_3_port, 
      Y_LOGIC_2_port, Y_LOGIC_1_port, Y_LOGIC_0_port, N111, N112, N113, 
      OUT_SHIFTER_31_port, OUT_SHIFTER_30_port, OUT_SHIFTER_29_port, 
      OUT_SHIFTER_28_port, OUT_SHIFTER_27_port, OUT_SHIFTER_26_port, 
      OUT_SHIFTER_25_port, OUT_SHIFTER_24_port, OUT_SHIFTER_23_port, 
      OUT_SHIFTER_22_port, OUT_SHIFTER_21_port, OUT_SHIFTER_20_port, 
      OUT_SHIFTER_19_port, OUT_SHIFTER_18_port, OUT_SHIFTER_17_port, 
      OUT_SHIFTER_16_port, OUT_SHIFTER_15_port, OUT_SHIFTER_14_port, 
      OUT_SHIFTER_13_port, OUT_SHIFTER_12_port, OUT_SHIFTER_11_port, 
      OUT_SHIFTER_10_port, OUT_SHIFTER_9_port, OUT_SHIFTER_8_port, 
      OUT_SHIFTER_7_port, OUT_SHIFTER_6_port, OUT_SHIFTER_5_port, 
      OUT_SHIFTER_4_port, OUT_SHIFTER_3_port, OUT_SHIFTER_2_port, 
      OUT_SHIFTER_1_port, OUT_SHIFTER_0_port, S_3_port, S_2_port, L0_31_port, 
      L0_30_port, L0_29_port, L0_28_port, L0_27_port, L0_26_port, L0_25_port, 
      L0_24_port, L0_23_port, L0_22_port, L0_21_port, L0_20_port, L0_19_port, 
      L0_18_port, L0_17_port, L0_16_port, L0_15_port, L0_14_port, L0_13_port, 
      L0_12_port, L0_11_port, L0_10_port, L0_9_port, L0_8_port, L0_7_port, 
      L0_6_port, L0_5_port, L0_4_port, L0_3_port, L0_2_port, L0_1_port, 
      L0_0_port, L1_31_port, L1_30_port, L1_29_port, L1_28_port, L1_27_port, 
      L1_26_port, L1_25_port, L1_24_port, L1_23_port, L1_22_port, L1_21_port, 
      L1_20_port, L1_19_port, L1_18_port, L1_17_port, L1_16_port, L1_15_port, 
      L1_14_port, L1_13_port, L1_12_port, L1_11_port, L1_10_port, L1_9_port, 
      L1_8_port, L1_7_port, L1_6_port, L1_5_port, L1_4_port, L1_3_port, 
      L1_2_port, L1_1_port, L1_0_port, L2_31_port, L2_30_port, L2_29_port, 
      L2_28_port, L2_27_port, L2_26_port, L2_25_port, L2_24_port, L2_23_port, 
      L2_22_port, L2_21_port, L2_20_port, L2_19_port, L2_18_port, L2_17_port, 
      L2_16_port, L2_15_port, L2_14_port, L2_13_port, L2_12_port, L2_11_port, 
      L2_10_port, L2_9_port, L2_8_port, L2_7_port, L2_6_port, L2_5_port, 
      L2_4_port, L2_3_port, L2_2_port, L2_1_port, L2_0_port, L3_31_port, 
      L3_30_port, L3_29_port, L3_28_port, L3_27_port, L3_26_port, L3_25_port, 
      L3_24_port, L3_23_port, L3_22_port, L3_21_port, L3_20_port, L3_19_port, 
      L3_18_port, L3_17_port, L3_16_port, L3_15_port, L3_14_port, L3_13_port, 
      L3_12_port, L3_11_port, L3_10_port, L3_9_port, L3_8_port, L3_7_port, 
      L3_6_port, L3_5_port, L3_4_port, L3_3_port, L3_2_port, L3_1_port, 
      L3_0_port, U2_U1_Z_0, U2_U2_Z_0, n12, n160, n1, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n84_port, n85_port, n86_port, n87_port, n88_port, n89_port, n90_port, 
      n91_port, n92_port, n93_port, n94_port, n95_port, n96_port, n97_port, 
      n98_port, n99_port, n100_port, n101_port, n102_port, n103_port, n104_port
      , n105_port, n106_port, n107_port, n108_port, n109_port, n110_port, 
      n111_port, n112_port, n113_port, n114, n115, n116, n117, n118, n119, n120
      , n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n_1050, n_1051, n_1052, n_1053 : std_logic;

begin
   
   X_Logic0_port <= '0';
   n12 <= '0';
   NAND31I_1 : NAND3_0 port map( A => n115, B => n147, C => X_Logic0_port, Y =>
                           L0_0_port);
   NAND31I_2 : NAND3_127 port map( A => n114, B => n146, C => X_Logic0_port, Y 
                           => L0_1_port);
   NAND31I_3 : NAND3_126 port map( A => n113_port, B => n145, C => 
                           X_Logic0_port, Y => L0_2_port);
   NAND31I_4 : NAND3_125 port map( A => n112_port, B => n144, C => 
                           X_Logic0_port, Y => L0_3_port);
   NAND31I_5 : NAND3_124 port map( A => n111_port, B => n143, C => 
                           X_Logic0_port, Y => L0_4_port);
   NAND31I_6 : NAND3_123 port map( A => n110_port, B => n142, C => 
                           X_Logic0_port, Y => L0_5_port);
   NAND31I_7 : NAND3_122 port map( A => n109_port, B => n141, C => 
                           X_Logic0_port, Y => L0_6_port);
   NAND31I_8 : NAND3_121 port map( A => n108_port, B => n140, C => 
                           X_Logic0_port, Y => L0_7_port);
   NAND31I_9 : NAND3_120 port map( A => n107_port, B => n139, C => 
                           X_Logic0_port, Y => L0_8_port);
   NAND31I_10 : NAND3_119 port map( A => n106_port, B => n138, C => 
                           X_Logic0_port, Y => L0_9_port);
   NAND31I_11 : NAND3_118 port map( A => n105_port, B => n137, C => 
                           X_Logic0_port, Y => L0_10_port);
   NAND31I_12 : NAND3_117 port map( A => n104_port, B => n136, C => 
                           X_Logic0_port, Y => L0_11_port);
   NAND31I_13 : NAND3_116 port map( A => n103_port, B => n135, C => 
                           X_Logic0_port, Y => L0_12_port);
   NAND31I_14 : NAND3_115 port map( A => n102_port, B => n134, C => 
                           X_Logic0_port, Y => L0_13_port);
   NAND31I_15 : NAND3_114 port map( A => n101_port, B => n133, C => 
                           X_Logic0_port, Y => L0_14_port);
   NAND31I_16 : NAND3_113 port map( A => n100_port, B => n132, C => 
                           X_Logic0_port, Y => L0_15_port);
   NAND31I_17 : NAND3_112 port map( A => n99_port, B => n131, C => 
                           X_Logic0_port, Y => L0_16_port);
   NAND31I_18 : NAND3_111 port map( A => n98_port, B => n130, C => 
                           X_Logic0_port, Y => L0_17_port);
   NAND31I_19 : NAND3_110 port map( A => n97_port, B => n129, C => 
                           X_Logic0_port, Y => L0_18_port);
   NAND31I_20 : NAND3_109 port map( A => n96_port, B => n128, C => 
                           X_Logic0_port, Y => L0_19_port);
   NAND31I_21 : NAND3_108 port map( A => n95_port, B => n127, C => 
                           X_Logic0_port, Y => L0_20_port);
   NAND31I_22 : NAND3_107 port map( A => n94_port, B => n126, C => 
                           X_Logic0_port, Y => L0_21_port);
   NAND31I_23 : NAND3_106 port map( A => n93_port, B => n125, C => 
                           X_Logic0_port, Y => L0_22_port);
   NAND31I_24 : NAND3_105 port map( A => n92_port, B => n124, C => 
                           X_Logic0_port, Y => L0_23_port);
   NAND31I_25 : NAND3_104 port map( A => n91_port, B => n123, C => 
                           X_Logic0_port, Y => L0_24_port);
   NAND31I_26 : NAND3_103 port map( A => n90_port, B => n122, C => 
                           X_Logic0_port, Y => L0_25_port);
   NAND31I_27 : NAND3_102 port map( A => n89_port, B => n121, C => 
                           X_Logic0_port, Y => L0_26_port);
   NAND31I_28 : NAND3_101 port map( A => n88_port, B => n120, C => 
                           X_Logic0_port, Y => L0_27_port);
   NAND31I_29 : NAND3_100 port map( A => n87_port, B => n119, C => 
                           X_Logic0_port, Y => L0_28_port);
   NAND31I_30 : NAND3_99 port map( A => n86_port, B => n118, C => X_Logic0_port
                           , Y => L0_29_port);
   NAND31I_31 : NAND3_98 port map( A => n85_port, B => n117, C => X_Logic0_port
                           , Y => L0_30_port);
   NAND31I_32 : NAND3_97 port map( A => n84_port, B => n116, C => X_Logic0_port
                           , Y => L0_31_port);
   NAND31I_1_0 : NAND3_96 port map( A => n115, B => DATA2(0), C => S_2_port, Y 
                           => L1_0_port);
   NAND31I_2_0 : NAND3_95 port map( A => n114, B => DATA2(1), C => S_2_port, Y 
                           => L1_1_port);
   NAND31I_3_0 : NAND3_94 port map( A => n113_port, B => DATA2(2), C => 
                           S_2_port, Y => L1_2_port);
   NAND31I_4_0 : NAND3_93 port map( A => n112_port, B => DATA2(3), C => 
                           S_2_port, Y => L1_3_port);
   NAND31I_5_0 : NAND3_92 port map( A => n111_port, B => DATA2(4), C => 
                           S_2_port, Y => L1_4_port);
   NAND31I_6_0 : NAND3_91 port map( A => n110_port, B => DATA2(5), C => 
                           S_2_port, Y => L1_5_port);
   NAND31I_7_0 : NAND3_90 port map( A => n109_port, B => DATA2(6), C => 
                           S_2_port, Y => L1_6_port);
   NAND31I_8_0 : NAND3_89 port map( A => n108_port, B => DATA2(7), C => 
                           S_2_port, Y => L1_7_port);
   NAND31I_9_0 : NAND3_88 port map( A => n107_port, B => DATA2(8), C => 
                           S_2_port, Y => L1_8_port);
   NAND31I_10_0 : NAND3_87 port map( A => n106_port, B => DATA2(9), C => 
                           S_2_port, Y => L1_9_port);
   NAND31I_11_0 : NAND3_86 port map( A => n105_port, B => DATA2(10), C => 
                           S_2_port, Y => L1_10_port);
   NAND31I_12_0 : NAND3_85 port map( A => n104_port, B => DATA2(11), C => 
                           S_2_port, Y => L1_11_port);
   NAND31I_13_0 : NAND3_84 port map( A => n103_port, B => DATA2(12), C => 
                           S_2_port, Y => L1_12_port);
   NAND31I_14_0 : NAND3_83 port map( A => n102_port, B => DATA2(13), C => 
                           S_2_port, Y => L1_13_port);
   NAND31I_15_0 : NAND3_82 port map( A => n101_port, B => DATA2(14), C => 
                           S_2_port, Y => L1_14_port);
   NAND31I_16_0 : NAND3_81 port map( A => n100_port, B => DATA2(15), C => 
                           S_2_port, Y => L1_15_port);
   NAND31I_17_0 : NAND3_80 port map( A => n99_port, B => DATA2(16), C => 
                           S_2_port, Y => L1_16_port);
   NAND31I_18_0 : NAND3_79 port map( A => n98_port, B => DATA2(17), C => 
                           S_2_port, Y => L1_17_port);
   NAND31I_19_0 : NAND3_78 port map( A => n97_port, B => DATA2(18), C => 
                           S_2_port, Y => L1_18_port);
   NAND31I_20_0 : NAND3_77 port map( A => n96_port, B => DATA2(19), C => 
                           S_2_port, Y => L1_19_port);
   NAND31I_21_0 : NAND3_76 port map( A => n95_port, B => DATA2(20), C => 
                           S_2_port, Y => L1_20_port);
   NAND31I_22_0 : NAND3_75 port map( A => n94_port, B => DATA2(21), C => 
                           S_2_port, Y => L1_21_port);
   NAND31I_23_0 : NAND3_74 port map( A => n93_port, B => DATA2(22), C => 
                           S_2_port, Y => L1_22_port);
   NAND31I_24_0 : NAND3_73 port map( A => n92_port, B => DATA2(23), C => 
                           S_2_port, Y => L1_23_port);
   NAND31I_25_0 : NAND3_72 port map( A => n91_port, B => DATA2(24), C => 
                           S_2_port, Y => L1_24_port);
   NAND31I_26_0 : NAND3_71 port map( A => n90_port, B => DATA2(25), C => 
                           S_2_port, Y => L1_25_port);
   NAND31I_27_0 : NAND3_70 port map( A => n89_port, B => DATA2(26), C => 
                           S_2_port, Y => L1_26_port);
   NAND31I_28_0 : NAND3_69 port map( A => n88_port, B => DATA2(27), C => 
                           S_2_port, Y => L1_27_port);
   NAND31I_29_0 : NAND3_68 port map( A => n87_port, B => DATA2(28), C => 
                           S_2_port, Y => L1_28_port);
   NAND31I_30_0 : NAND3_67 port map( A => n86_port, B => DATA2(29), C => 
                           S_2_port, Y => L1_29_port);
   NAND31I_31_0 : NAND3_66 port map( A => n85_port, B => DATA2(30), C => 
                           S_2_port, Y => L1_30_port);
   NAND31I_32_0 : NAND3_65 port map( A => n84_port, B => DATA2(31), C => 
                           S_2_port, Y => L1_31_port);
   NAND31I_1_1 : NAND3_64 port map( A => DATA1(0), B => n147, C => S_2_port, Y 
                           => L2_0_port);
   NAND31I_2_1 : NAND3_63 port map( A => DATA1(1), B => n146, C => S_2_port, Y 
                           => L2_1_port);
   NAND31I_3_1 : NAND3_62 port map( A => DATA1(2), B => n145, C => S_2_port, Y 
                           => L2_2_port);
   NAND31I_4_1 : NAND3_61 port map( A => DATA1(3), B => n144, C => S_2_port, Y 
                           => L2_3_port);
   NAND31I_5_1 : NAND3_60 port map( A => DATA1(4), B => n143, C => S_2_port, Y 
                           => L2_4_port);
   NAND31I_6_1 : NAND3_59 port map( A => DATA1(5), B => n142, C => S_2_port, Y 
                           => L2_5_port);
   NAND31I_7_1 : NAND3_58 port map( A => DATA1(6), B => n141, C => S_2_port, Y 
                           => L2_6_port);
   NAND31I_8_1 : NAND3_57 port map( A => DATA1(7), B => n140, C => S_2_port, Y 
                           => L2_7_port);
   NAND31I_9_1 : NAND3_56 port map( A => DATA1(8), B => n139, C => S_2_port, Y 
                           => L2_8_port);
   NAND31I_10_1 : NAND3_55 port map( A => DATA1(9), B => n138, C => S_2_port, Y
                           => L2_9_port);
   NAND31I_11_1 : NAND3_54 port map( A => DATA1(10), B => n137, C => S_2_port, 
                           Y => L2_10_port);
   NAND31I_12_1 : NAND3_53 port map( A => DATA1(11), B => n136, C => S_2_port, 
                           Y => L2_11_port);
   NAND31I_13_1 : NAND3_52 port map( A => DATA1(12), B => n135, C => S_2_port, 
                           Y => L2_12_port);
   NAND31I_14_1 : NAND3_51 port map( A => DATA1(13), B => n134, C => S_2_port, 
                           Y => L2_13_port);
   NAND31I_15_1 : NAND3_50 port map( A => DATA1(14), B => n133, C => S_2_port, 
                           Y => L2_14_port);
   NAND31I_16_1 : NAND3_49 port map( A => DATA1(15), B => n132, C => S_2_port, 
                           Y => L2_15_port);
   NAND31I_17_1 : NAND3_48 port map( A => DATA1(16), B => n131, C => S_2_port, 
                           Y => L2_16_port);
   NAND31I_18_1 : NAND3_47 port map( A => DATA1(17), B => n130, C => S_2_port, 
                           Y => L2_17_port);
   NAND31I_19_1 : NAND3_46 port map( A => DATA1(18), B => n129, C => S_2_port, 
                           Y => L2_18_port);
   NAND31I_20_1 : NAND3_45 port map( A => DATA1(19), B => n128, C => S_2_port, 
                           Y => L2_19_port);
   NAND31I_21_1 : NAND3_44 port map( A => DATA1(20), B => n127, C => S_2_port, 
                           Y => L2_20_port);
   NAND31I_22_1 : NAND3_43 port map( A => DATA1(21), B => n126, C => S_2_port, 
                           Y => L2_21_port);
   NAND31I_23_1 : NAND3_42 port map( A => DATA1(22), B => n125, C => S_2_port, 
                           Y => L2_22_port);
   NAND31I_24_1 : NAND3_41 port map( A => DATA1(23), B => n124, C => S_2_port, 
                           Y => L2_23_port);
   NAND31I_25_1 : NAND3_40 port map( A => DATA1(24), B => n123, C => S_2_port, 
                           Y => L2_24_port);
   NAND31I_26_1 : NAND3_39 port map( A => DATA1(25), B => n122, C => S_2_port, 
                           Y => L2_25_port);
   NAND31I_27_1 : NAND3_38 port map( A => DATA1(26), B => n121, C => S_2_port, 
                           Y => L2_26_port);
   NAND31I_28_1 : NAND3_37 port map( A => DATA1(27), B => n120, C => S_2_port, 
                           Y => L2_27_port);
   NAND31I_29_1 : NAND3_36 port map( A => DATA1(28), B => n119, C => S_2_port, 
                           Y => L2_28_port);
   NAND31I_30_1 : NAND3_35 port map( A => DATA1(29), B => n118, C => S_2_port, 
                           Y => L2_29_port);
   NAND31I_31_1 : NAND3_34 port map( A => DATA1(30), B => n117, C => S_2_port, 
                           Y => L2_30_port);
   NAND31I_32_1 : NAND3_33 port map( A => DATA1(31), B => n116, C => S_2_port, 
                           Y => L2_31_port);
   NAND31I_1_2 : NAND3_32 port map( A => DATA1(0), B => DATA2(0), C => S_3_port
                           , Y => L3_0_port);
   NAND31I_2_2 : NAND3_31 port map( A => DATA1(1), B => DATA2(1), C => S_3_port
                           , Y => L3_1_port);
   NAND31I_3_2 : NAND3_30 port map( A => DATA1(2), B => DATA2(2), C => S_3_port
                           , Y => L3_2_port);
   NAND31I_4_2 : NAND3_29 port map( A => DATA1(3), B => DATA2(3), C => S_3_port
                           , Y => L3_3_port);
   NAND31I_5_2 : NAND3_28 port map( A => DATA1(4), B => DATA2(4), C => S_3_port
                           , Y => L3_4_port);
   NAND31I_6_2 : NAND3_27 port map( A => DATA1(5), B => DATA2(5), C => S_3_port
                           , Y => L3_5_port);
   NAND31I_7_2 : NAND3_26 port map( A => DATA1(6), B => DATA2(6), C => S_3_port
                           , Y => L3_6_port);
   NAND31I_8_2 : NAND3_25 port map( A => DATA1(7), B => DATA2(7), C => S_3_port
                           , Y => L3_7_port);
   NAND31I_9_2 : NAND3_24 port map( A => DATA1(8), B => DATA2(8), C => S_3_port
                           , Y => L3_8_port);
   NAND31I_10_2 : NAND3_23 port map( A => DATA1(9), B => DATA2(9), C => 
                           S_3_port, Y => L3_9_port);
   NAND31I_11_2 : NAND3_22 port map( A => DATA1(10), B => DATA2(10), C => 
                           S_3_port, Y => L3_10_port);
   NAND31I_12_2 : NAND3_21 port map( A => DATA1(11), B => DATA2(11), C => 
                           S_3_port, Y => L3_11_port);
   NAND31I_13_2 : NAND3_20 port map( A => DATA1(12), B => DATA2(12), C => 
                           S_3_port, Y => L3_12_port);
   NAND31I_14_2 : NAND3_19 port map( A => DATA1(13), B => DATA2(13), C => 
                           S_3_port, Y => L3_13_port);
   NAND31I_15_2 : NAND3_18 port map( A => DATA1(14), B => DATA2(14), C => 
                           S_3_port, Y => L3_14_port);
   NAND31I_16_2 : NAND3_17 port map( A => DATA1(15), B => DATA2(15), C => 
                           S_3_port, Y => L3_15_port);
   NAND31I_17_2 : NAND3_16 port map( A => DATA1(16), B => DATA2(16), C => 
                           S_3_port, Y => L3_16_port);
   NAND31I_18_2 : NAND3_15 port map( A => DATA1(17), B => DATA2(17), C => 
                           S_3_port, Y => L3_17_port);
   NAND31I_19_2 : NAND3_14 port map( A => DATA1(18), B => DATA2(18), C => 
                           S_3_port, Y => L3_18_port);
   NAND31I_20_2 : NAND3_13 port map( A => DATA1(19), B => DATA2(19), C => 
                           S_3_port, Y => L3_19_port);
   NAND31I_21_2 : NAND3_12 port map( A => DATA1(20), B => DATA2(20), C => 
                           S_3_port, Y => L3_20_port);
   NAND31I_22_2 : NAND3_11 port map( A => DATA1(21), B => DATA2(21), C => 
                           S_3_port, Y => L3_21_port);
   NAND31I_23_2 : NAND3_10 port map( A => DATA1(22), B => DATA2(22), C => 
                           S_3_port, Y => L3_22_port);
   NAND31I_24_2 : NAND3_9 port map( A => DATA1(23), B => DATA2(23), C => 
                           S_3_port, Y => L3_23_port);
   NAND31I_25_2 : NAND3_8 port map( A => DATA1(24), B => DATA2(24), C => 
                           S_3_port, Y => L3_24_port);
   NAND31I_26_2 : NAND3_7 port map( A => DATA1(25), B => DATA2(25), C => 
                           S_3_port, Y => L3_25_port);
   NAND31I_27_2 : NAND3_6 port map( A => DATA1(26), B => DATA2(26), C => 
                           S_3_port, Y => L3_26_port);
   NAND31I_28_2 : NAND3_5 port map( A => DATA1(27), B => DATA2(27), C => 
                           S_3_port, Y => L3_27_port);
   NAND31I_29_2 : NAND3_4 port map( A => DATA1(28), B => DATA2(28), C => 
                           S_3_port, Y => L3_28_port);
   NAND31I_30_2 : NAND3_3 port map( A => DATA1(29), B => DATA2(29), C => 
                           S_3_port, Y => L3_29_port);
   NAND31I_31_2 : NAND3_2 port map( A => DATA1(30), B => DATA2(30), C => 
                           S_3_port, Y => L3_30_port);
   NAND31I_32_2 : NAND3_1 port map( A => DATA1(31), B => DATA2(31), C => 
                           S_3_port, Y => L3_31_port);
   NAND41I_1 : NAND4_0 port map( A => L0_0_port, B => L1_0_port, C => L2_0_port
                           , D => L3_0_port, Y => Y_LOGIC_0_port);
   NAND41I_2 : NAND4_31 port map( A => L0_1_port, B => L1_1_port, C => 
                           L2_1_port, D => L3_1_port, Y => Y_LOGIC_1_port);
   NAND41I_3 : NAND4_30 port map( A => L0_2_port, B => L1_2_port, C => 
                           L2_2_port, D => L3_2_port, Y => Y_LOGIC_2_port);
   NAND41I_4 : NAND4_29 port map( A => L0_3_port, B => L1_3_port, C => 
                           L2_3_port, D => L3_3_port, Y => Y_LOGIC_3_port);
   NAND41I_5 : NAND4_28 port map( A => L0_4_port, B => L1_4_port, C => 
                           L2_4_port, D => L3_4_port, Y => Y_LOGIC_4_port);
   NAND41I_6 : NAND4_27 port map( A => L0_5_port, B => L1_5_port, C => 
                           L2_5_port, D => L3_5_port, Y => Y_LOGIC_5_port);
   NAND41I_7 : NAND4_26 port map( A => L0_6_port, B => L1_6_port, C => 
                           L2_6_port, D => L3_6_port, Y => Y_LOGIC_6_port);
   NAND41I_8 : NAND4_25 port map( A => L0_7_port, B => L1_7_port, C => 
                           L2_7_port, D => L3_7_port, Y => Y_LOGIC_7_port);
   NAND41I_9 : NAND4_24 port map( A => L0_8_port, B => L1_8_port, C => 
                           L2_8_port, D => L3_8_port, Y => Y_LOGIC_8_port);
   NAND41I_10 : NAND4_23 port map( A => L0_9_port, B => L1_9_port, C => 
                           L2_9_port, D => L3_9_port, Y => Y_LOGIC_9_port);
   NAND41I_11 : NAND4_22 port map( A => L0_10_port, B => L1_10_port, C => 
                           L2_10_port, D => L3_10_port, Y => Y_LOGIC_10_port);
   NAND41I_12 : NAND4_21 port map( A => L0_11_port, B => L1_11_port, C => 
                           L2_11_port, D => L3_11_port, Y => Y_LOGIC_11_port);
   NAND41I_13 : NAND4_20 port map( A => L0_12_port, B => L1_12_port, C => 
                           L2_12_port, D => L3_12_port, Y => Y_LOGIC_12_port);
   NAND41I_14 : NAND4_19 port map( A => L0_13_port, B => L1_13_port, C => 
                           L2_13_port, D => L3_13_port, Y => Y_LOGIC_13_port);
   NAND41I_15 : NAND4_18 port map( A => L0_14_port, B => L1_14_port, C => 
                           L2_14_port, D => L3_14_port, Y => Y_LOGIC_14_port);
   NAND41I_16 : NAND4_17 port map( A => L0_15_port, B => L1_15_port, C => 
                           L2_15_port, D => L3_15_port, Y => Y_LOGIC_15_port);
   NAND41I_17 : NAND4_16 port map( A => L0_16_port, B => L1_16_port, C => 
                           L2_16_port, D => L3_16_port, Y => Y_LOGIC_16_port);
   NAND41I_18 : NAND4_15 port map( A => L0_17_port, B => L1_17_port, C => 
                           L2_17_port, D => L3_17_port, Y => Y_LOGIC_17_port);
   NAND41I_19 : NAND4_14 port map( A => L0_18_port, B => L1_18_port, C => 
                           L2_18_port, D => L3_18_port, Y => Y_LOGIC_18_port);
   NAND41I_20 : NAND4_13 port map( A => L0_19_port, B => L1_19_port, C => 
                           L2_19_port, D => L3_19_port, Y => Y_LOGIC_19_port);
   NAND41I_21 : NAND4_12 port map( A => L0_20_port, B => L1_20_port, C => 
                           L2_20_port, D => L3_20_port, Y => Y_LOGIC_20_port);
   NAND41I_22 : NAND4_11 port map( A => L0_21_port, B => L1_21_port, C => 
                           L2_21_port, D => L3_21_port, Y => Y_LOGIC_21_port);
   NAND41I_23 : NAND4_10 port map( A => L0_22_port, B => L1_22_port, C => 
                           L2_22_port, D => L3_22_port, Y => Y_LOGIC_22_port);
   NAND41I_24 : NAND4_9 port map( A => L0_23_port, B => L1_23_port, C => 
                           L2_23_port, D => L3_23_port, Y => Y_LOGIC_23_port);
   NAND41I_25 : NAND4_8 port map( A => L0_24_port, B => L1_24_port, C => 
                           L2_24_port, D => L3_24_port, Y => Y_LOGIC_24_port);
   NAND41I_26 : NAND4_7 port map( A => L0_25_port, B => L1_25_port, C => 
                           L2_25_port, D => L3_25_port, Y => Y_LOGIC_25_port);
   NAND41I_27 : NAND4_6 port map( A => L0_26_port, B => L1_26_port, C => 
                           L2_26_port, D => L3_26_port, Y => Y_LOGIC_26_port);
   NAND41I_28 : NAND4_5 port map( A => L0_27_port, B => L1_27_port, C => 
                           L2_27_port, D => L3_27_port, Y => Y_LOGIC_27_port);
   NAND41I_29 : NAND4_4 port map( A => L0_28_port, B => L1_28_port, C => 
                           L2_28_port, D => L3_28_port, Y => Y_LOGIC_28_port);
   NAND41I_30 : NAND4_3 port map( A => L0_29_port, B => L1_29_port, C => 
                           L2_29_port, D => L3_29_port, Y => Y_LOGIC_29_port);
   NAND41I_31 : NAND4_2 port map( A => L0_30_port, B => L1_30_port, C => 
                           L2_30_port, D => L3_30_port, Y => Y_LOGIC_30_port);
   NAND41I_32 : NAND4_1 port map( A => L0_31_port, B => L1_31_port, C => 
                           L2_31_port, D => L3_31_port, Y => Y_LOGIC_31_port);
   SHIFTER : BARREL_SHIFTER_N32 port map( CONF => n160, DATA1(31) => DATA1(31),
                           DATA1(30) => DATA1(30), DATA1(29) => DATA1(29), 
                           DATA1(28) => DATA1(28), DATA1(27) => DATA1(27), 
                           DATA1(26) => DATA1(26), DATA1(25) => DATA1(25), 
                           DATA1(24) => DATA1(24), DATA1(23) => DATA1(23), 
                           DATA1(22) => DATA1(22), DATA1(21) => DATA1(21), 
                           DATA1(20) => DATA1(20), DATA1(19) => DATA1(19), 
                           DATA1(18) => DATA1(18), DATA1(17) => DATA1(17), 
                           DATA1(16) => DATA1(16), DATA1(15) => DATA1(15), 
                           DATA1(14) => DATA1(14), DATA1(13) => DATA1(13), 
                           DATA1(12) => DATA1(12), DATA1(11) => DATA1(11), 
                           DATA1(10) => DATA1(10), DATA1(9) => DATA1(9), 
                           DATA1(8) => DATA1(8), DATA1(7) => DATA1(7), DATA1(6)
                           => DATA1(6), DATA1(5) => DATA1(5), DATA1(4) => 
                           DATA1(4), DATA1(3) => DATA1(3), DATA1(2) => DATA1(2)
                           , DATA1(1) => DATA1(1), DATA1(0) => DATA1(0), 
                           DATA2(31) => DATA2(31), DATA2(30) => DATA2(30), 
                           DATA2(29) => DATA2(29), DATA2(28) => DATA2(28), 
                           DATA2(27) => DATA2(27), DATA2(26) => DATA2(26), 
                           DATA2(25) => DATA2(25), DATA2(24) => DATA2(24), 
                           DATA2(23) => DATA2(23), DATA2(22) => DATA2(22), 
                           DATA2(21) => DATA2(21), DATA2(20) => DATA2(20), 
                           DATA2(19) => DATA2(19), DATA2(18) => DATA2(18), 
                           DATA2(17) => DATA2(17), DATA2(16) => DATA2(16), 
                           DATA2(15) => DATA2(15), DATA2(14) => DATA2(14), 
                           DATA2(13) => DATA2(13), DATA2(12) => DATA2(12), 
                           DATA2(11) => DATA2(11), DATA2(10) => DATA2(10), 
                           DATA2(9) => DATA2(9), DATA2(8) => DATA2(8), DATA2(7)
                           => DATA2(7), DATA2(6) => DATA2(6), DATA2(5) => 
                           DATA2(5), DATA2(4) => DATA2(4), DATA2(3) => DATA2(3)
                           , DATA2(2) => DATA2(2), DATA2(1) => DATA2(1), 
                           DATA2(0) => DATA2(0), OUTPUT(31) => 
                           OUT_SHIFTER_31_port, OUTPUT(30) => 
                           OUT_SHIFTER_30_port, OUTPUT(29) => 
                           OUT_SHIFTER_29_port, OUTPUT(28) => 
                           OUT_SHIFTER_28_port, OUTPUT(27) => 
                           OUT_SHIFTER_27_port, OUTPUT(26) => 
                           OUT_SHIFTER_26_port, OUTPUT(25) => 
                           OUT_SHIFTER_25_port, OUTPUT(24) => 
                           OUT_SHIFTER_24_port, OUTPUT(23) => 
                           OUT_SHIFTER_23_port, OUTPUT(22) => 
                           OUT_SHIFTER_22_port, OUTPUT(21) => 
                           OUT_SHIFTER_21_port, OUTPUT(20) => 
                           OUT_SHIFTER_20_port, OUTPUT(19) => 
                           OUT_SHIFTER_19_port, OUTPUT(18) => 
                           OUT_SHIFTER_18_port, OUTPUT(17) => 
                           OUT_SHIFTER_17_port, OUTPUT(16) => 
                           OUT_SHIFTER_16_port, OUTPUT(15) => 
                           OUT_SHIFTER_15_port, OUTPUT(14) => 
                           OUT_SHIFTER_14_port, OUTPUT(13) => 
                           OUT_SHIFTER_13_port, OUTPUT(12) => 
                           OUT_SHIFTER_12_port, OUTPUT(11) => 
                           OUT_SHIFTER_11_port, OUTPUT(10) => 
                           OUT_SHIFTER_10_port, OUTPUT(9) => OUT_SHIFTER_9_port
                           , OUTPUT(8) => OUT_SHIFTER_8_port, OUTPUT(7) => 
                           OUT_SHIFTER_7_port, OUTPUT(6) => OUT_SHIFTER_6_port,
                           OUTPUT(5) => OUT_SHIFTER_5_port, OUTPUT(4) => 
                           OUT_SHIFTER_4_port, OUTPUT(3) => OUT_SHIFTER_3_port,
                           OUTPUT(2) => OUT_SHIFTER_2_port, OUTPUT(1) => 
                           OUT_SHIFTER_1_port, OUTPUT(0) => OUT_SHIFTER_0_port)
                           ;
   r75 : ALU_N32_DW01_addsub_0 port map( A(31) => DATA1(31), A(30) => DATA1(30)
                           , A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , CI => n12, ADD_SUB => U2_U1_Z_0, SUM(31) => N110, 
                           SUM(30) => N109, SUM(29) => N108, SUM(28) => N107, 
                           SUM(27) => N106, SUM(26) => N105, SUM(25) => N104, 
                           SUM(24) => N103, SUM(23) => N102, SUM(22) => N101, 
                           SUM(21) => N100, SUM(20) => N99, SUM(19) => N98, 
                           SUM(18) => N97, SUM(17) => N96, SUM(16) => N95, 
                           SUM(15) => N94, SUM(14) => N93, SUM(13) => N92, 
                           SUM(12) => N91, SUM(11) => N90, SUM(10) => N89, 
                           SUM(9) => N88, SUM(8) => N87, SUM(7) => N86, SUM(6) 
                           => N85, SUM(5) => N84, SUM(4) => N83, SUM(3) => N82,
                           SUM(2) => N81, SUM(1) => N80, SUM(0) => N79, CO => 
                           n_1050);
   r69 : ALU_N32_DW01_cmp6_0 port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , TC => U2_U2_Z_0, LT => n_1051, GT => n_1052, EQ =>
                           n_1053, LE => N111, GE => N112, NE => N113);
   U3 : INV_X4 port map( A => n38, ZN => S_2_port);
   U4 : NAND2_X2 port map( A1 => n38, A2 => n39, ZN => n4);
   U5 : NAND2_X2 port map( A1 => n37, A2 => n46, ZN => n3);
   U6 : NAND2_X2 port map( A1 => n36, A2 => n48, ZN => n2);
   U7 : INV_X2 port map( A => n37, ZN => U2_U1_Z_0);
   U8 : OAI21_X4 port map( B1 => FUNC(3), B2 => n38, A => n39, ZN => S_3_port);
   U9 : INV_X1 port map( A => n1, ZN => OUTALU(31));
   U10 : AOI222_X1 port map( A1 => OUT_SHIFTER_31_port, A2 => n2, B1 => N110, 
                           B2 => n3, C1 => Y_LOGIC_31_port, C2 => n4, ZN => n1)
                           ;
   U11 : INV_X1 port map( A => n5, ZN => OUTALU(30));
   U12 : AOI222_X1 port map( A1 => OUT_SHIFTER_30_port, A2 => n2, B1 => N109, 
                           B2 => n3, C1 => Y_LOGIC_30_port, C2 => n4, ZN => n5)
                           ;
   U13 : INV_X1 port map( A => n6, ZN => OUTALU(29));
   U14 : AOI222_X1 port map( A1 => OUT_SHIFTER_29_port, A2 => n2, B1 => N108, 
                           B2 => n3, C1 => Y_LOGIC_29_port, C2 => n4, ZN => n6)
                           ;
   U15 : INV_X1 port map( A => n7, ZN => OUTALU(28));
   U16 : AOI222_X1 port map( A1 => OUT_SHIFTER_28_port, A2 => n2, B1 => N107, 
                           B2 => n3, C1 => Y_LOGIC_28_port, C2 => n4, ZN => n7)
                           ;
   U17 : INV_X1 port map( A => n8, ZN => OUTALU(27));
   U18 : AOI222_X1 port map( A1 => OUT_SHIFTER_27_port, A2 => n2, B1 => N106, 
                           B2 => n3, C1 => Y_LOGIC_27_port, C2 => n4, ZN => n8)
                           ;
   U19 : INV_X1 port map( A => n9, ZN => OUTALU(26));
   U20 : AOI222_X1 port map( A1 => OUT_SHIFTER_26_port, A2 => n2, B1 => N105, 
                           B2 => n3, C1 => Y_LOGIC_26_port, C2 => n4, ZN => n9)
                           ;
   U21 : INV_X1 port map( A => n10, ZN => OUTALU(25));
   U22 : AOI222_X1 port map( A1 => OUT_SHIFTER_25_port, A2 => n2, B1 => N104, 
                           B2 => n3, C1 => Y_LOGIC_25_port, C2 => n4, ZN => n10
                           );
   U23 : INV_X1 port map( A => n11, ZN => OUTALU(24));
   U24 : AOI222_X1 port map( A1 => OUT_SHIFTER_24_port, A2 => n2, B1 => N103, 
                           B2 => n3, C1 => Y_LOGIC_24_port, C2 => n4, ZN => n11
                           );
   U25 : INV_X1 port map( A => n13, ZN => OUTALU(23));
   U26 : AOI222_X1 port map( A1 => OUT_SHIFTER_23_port, A2 => n2, B1 => N102, 
                           B2 => n3, C1 => Y_LOGIC_23_port, C2 => n4, ZN => n13
                           );
   U27 : INV_X1 port map( A => n14, ZN => OUTALU(14));
   U28 : AOI222_X1 port map( A1 => OUT_SHIFTER_14_port, A2 => n2, B1 => N93, B2
                           => n3, C1 => Y_LOGIC_14_port, C2 => n4, ZN => n14);
   U29 : INV_X1 port map( A => n15, ZN => OUTALU(13));
   U30 : AOI222_X1 port map( A1 => OUT_SHIFTER_13_port, A2 => n2, B1 => N92, B2
                           => n3, C1 => Y_LOGIC_13_port, C2 => n4, ZN => n15);
   U31 : INV_X1 port map( A => n16, ZN => OUTALU(12));
   U32 : AOI222_X1 port map( A1 => OUT_SHIFTER_12_port, A2 => n2, B1 => N91, B2
                           => n3, C1 => Y_LOGIC_12_port, C2 => n4, ZN => n16);
   U33 : INV_X1 port map( A => n17, ZN => OUTALU(11));
   U34 : AOI222_X1 port map( A1 => OUT_SHIFTER_11_port, A2 => n2, B1 => N90, B2
                           => n3, C1 => Y_LOGIC_11_port, C2 => n4, ZN => n17);
   U35 : INV_X1 port map( A => n18, ZN => OUTALU(10));
   U36 : AOI222_X1 port map( A1 => OUT_SHIFTER_10_port, A2 => n2, B1 => N89, B2
                           => n3, C1 => Y_LOGIC_10_port, C2 => n4, ZN => n18);
   U37 : INV_X1 port map( A => n19, ZN => OUTALU(9));
   U38 : AOI222_X1 port map( A1 => OUT_SHIFTER_9_port, A2 => n2, B1 => N88, B2 
                           => n3, C1 => Y_LOGIC_9_port, C2 => n4, ZN => n19);
   U39 : INV_X1 port map( A => n20, ZN => OUTALU(8));
   U40 : AOI222_X1 port map( A1 => OUT_SHIFTER_8_port, A2 => n2, B1 => N87, B2 
                           => n3, C1 => Y_LOGIC_8_port, C2 => n4, ZN => n20);
   U41 : INV_X1 port map( A => n21, ZN => OUTALU(7));
   U42 : AOI222_X1 port map( A1 => OUT_SHIFTER_7_port, A2 => n2, B1 => N86, B2 
                           => n3, C1 => Y_LOGIC_7_port, C2 => n4, ZN => n21);
   U43 : INV_X1 port map( A => n22, ZN => OUTALU(15));
   U44 : AOI222_X1 port map( A1 => OUT_SHIFTER_15_port, A2 => n2, B1 => N94, B2
                           => n3, C1 => Y_LOGIC_15_port, C2 => n4, ZN => n22);
   U45 : INV_X1 port map( A => n23, ZN => OUTALU(22));
   U46 : AOI222_X1 port map( A1 => OUT_SHIFTER_22_port, A2 => n2, B1 => N101, 
                           B2 => n3, C1 => Y_LOGIC_22_port, C2 => n4, ZN => n23
                           );
   U47 : INV_X1 port map( A => n24, ZN => OUTALU(21));
   U48 : AOI222_X1 port map( A1 => OUT_SHIFTER_21_port, A2 => n2, B1 => N100, 
                           B2 => n3, C1 => Y_LOGIC_21_port, C2 => n4, ZN => n24
                           );
   U49 : INV_X1 port map( A => n25, ZN => OUTALU(20));
   U50 : AOI222_X1 port map( A1 => OUT_SHIFTER_20_port, A2 => n2, B1 => N99, B2
                           => n3, C1 => Y_LOGIC_20_port, C2 => n4, ZN => n25);
   U51 : INV_X1 port map( A => n26, ZN => OUTALU(19));
   U52 : AOI222_X1 port map( A1 => OUT_SHIFTER_19_port, A2 => n2, B1 => N98, B2
                           => n3, C1 => Y_LOGIC_19_port, C2 => n4, ZN => n26);
   U53 : INV_X1 port map( A => n27, ZN => OUTALU(18));
   U54 : AOI222_X1 port map( A1 => OUT_SHIFTER_18_port, A2 => n2, B1 => N97, B2
                           => n3, C1 => Y_LOGIC_18_port, C2 => n4, ZN => n27);
   U55 : INV_X1 port map( A => n28, ZN => OUTALU(17));
   U56 : AOI222_X1 port map( A1 => OUT_SHIFTER_17_port, A2 => n2, B1 => N96, B2
                           => n3, C1 => Y_LOGIC_17_port, C2 => n4, ZN => n28);
   U57 : INV_X1 port map( A => n29, ZN => OUTALU(16));
   U58 : AOI222_X1 port map( A1 => OUT_SHIFTER_16_port, A2 => n2, B1 => N95, B2
                           => n3, C1 => Y_LOGIC_16_port, C2 => n4, ZN => n29);
   U59 : INV_X1 port map( A => n30, ZN => OUTALU(6));
   U60 : AOI222_X1 port map( A1 => OUT_SHIFTER_6_port, A2 => n2, B1 => N85, B2 
                           => n3, C1 => Y_LOGIC_6_port, C2 => n4, ZN => n30);
   U61 : INV_X1 port map( A => n31, ZN => OUTALU(5));
   U62 : AOI222_X1 port map( A1 => OUT_SHIFTER_5_port, A2 => n2, B1 => N84, B2 
                           => n3, C1 => Y_LOGIC_5_port, C2 => n4, ZN => n31);
   U63 : INV_X1 port map( A => n32, ZN => OUTALU(4));
   U64 : AOI222_X1 port map( A1 => OUT_SHIFTER_4_port, A2 => n2, B1 => N83, B2 
                           => n3, C1 => Y_LOGIC_4_port, C2 => n4, ZN => n32);
   U65 : INV_X1 port map( A => n33, ZN => OUTALU(3));
   U66 : AOI222_X1 port map( A1 => OUT_SHIFTER_3_port, A2 => n2, B1 => N82, B2 
                           => n3, C1 => Y_LOGIC_3_port, C2 => n4, ZN => n33);
   U67 : INV_X1 port map( A => n34, ZN => OUTALU(2));
   U68 : AOI222_X1 port map( A1 => OUT_SHIFTER_2_port, A2 => n2, B1 => N81, B2 
                           => n3, C1 => Y_LOGIC_2_port, C2 => n4, ZN => n34);
   U69 : INV_X1 port map( A => n35, ZN => OUTALU(1));
   U70 : AOI222_X1 port map( A1 => OUT_SHIFTER_1_port, A2 => n2, B1 => N80, B2 
                           => n3, C1 => Y_LOGIC_1_port, C2 => n4, ZN => n35);
   U71 : INV_X1 port map( A => DATA1(31), ZN => n84_port);
   U72 : INV_X1 port map( A => DATA1(30), ZN => n85_port);
   U73 : INV_X1 port map( A => DATA1(29), ZN => n86_port);
   U74 : INV_X1 port map( A => DATA1(28), ZN => n87_port);
   U75 : INV_X1 port map( A => DATA1(27), ZN => n88_port);
   U76 : INV_X1 port map( A => DATA1(26), ZN => n89_port);
   U77 : INV_X1 port map( A => DATA1(25), ZN => n90_port);
   U78 : INV_X1 port map( A => DATA1(24), ZN => n91_port);
   U79 : INV_X1 port map( A => DATA1(23), ZN => n92_port);
   U80 : INV_X1 port map( A => DATA1(22), ZN => n93_port);
   U81 : INV_X1 port map( A => DATA1(21), ZN => n94_port);
   U82 : INV_X1 port map( A => DATA1(20), ZN => n95_port);
   U83 : INV_X1 port map( A => DATA1(19), ZN => n96_port);
   U84 : INV_X1 port map( A => DATA1(18), ZN => n97_port);
   U85 : INV_X1 port map( A => DATA1(17), ZN => n98_port);
   U86 : INV_X1 port map( A => DATA1(16), ZN => n99_port);
   U87 : INV_X1 port map( A => DATA1(15), ZN => n100_port);
   U88 : INV_X1 port map( A => DATA1(14), ZN => n101_port);
   U89 : INV_X1 port map( A => DATA1(13), ZN => n102_port);
   U90 : INV_X1 port map( A => DATA1(12), ZN => n103_port);
   U91 : INV_X1 port map( A => DATA1(11), ZN => n104_port);
   U92 : INV_X1 port map( A => DATA1(10), ZN => n105_port);
   U93 : INV_X1 port map( A => DATA1(9), ZN => n106_port);
   U94 : INV_X1 port map( A => DATA1(8), ZN => n107_port);
   U95 : INV_X1 port map( A => DATA1(7), ZN => n108_port);
   U96 : INV_X1 port map( A => DATA1(6), ZN => n109_port);
   U97 : INV_X1 port map( A => DATA1(5), ZN => n110_port);
   U98 : INV_X1 port map( A => DATA1(4), ZN => n111_port);
   U99 : INV_X1 port map( A => DATA1(3), ZN => n112_port);
   U100 : INV_X1 port map( A => DATA1(2), ZN => n113_port);
   U101 : INV_X1 port map( A => DATA1(1), ZN => n114);
   U102 : INV_X1 port map( A => DATA1(0), ZN => n115);
   U103 : INV_X1 port map( A => DATA2(31), ZN => n116);
   U104 : INV_X1 port map( A => DATA2(30), ZN => n117);
   U105 : INV_X1 port map( A => DATA2(29), ZN => n118);
   U106 : INV_X1 port map( A => DATA2(28), ZN => n119);
   U107 : INV_X1 port map( A => DATA2(27), ZN => n120);
   U108 : INV_X1 port map( A => DATA2(26), ZN => n121);
   U109 : INV_X1 port map( A => DATA2(25), ZN => n122);
   U110 : INV_X1 port map( A => DATA2(24), ZN => n123);
   U111 : INV_X1 port map( A => DATA2(23), ZN => n124);
   U112 : INV_X1 port map( A => DATA2(22), ZN => n125);
   U113 : INV_X1 port map( A => DATA2(21), ZN => n126);
   U114 : INV_X1 port map( A => DATA2(20), ZN => n127);
   U115 : INV_X1 port map( A => DATA2(19), ZN => n128);
   U116 : INV_X1 port map( A => DATA2(18), ZN => n129);
   U117 : INV_X1 port map( A => DATA2(17), ZN => n130);
   U118 : INV_X1 port map( A => DATA2(16), ZN => n131);
   U119 : INV_X1 port map( A => DATA2(15), ZN => n132);
   U120 : INV_X1 port map( A => DATA2(14), ZN => n133);
   U121 : INV_X1 port map( A => DATA2(13), ZN => n134);
   U122 : INV_X1 port map( A => DATA2(12), ZN => n135);
   U123 : INV_X1 port map( A => DATA2(11), ZN => n136);
   U124 : INV_X1 port map( A => DATA2(10), ZN => n137);
   U125 : INV_X1 port map( A => DATA2(9), ZN => n138);
   U126 : INV_X1 port map( A => DATA2(8), ZN => n139);
   U127 : INV_X1 port map( A => DATA2(7), ZN => n140);
   U128 : INV_X1 port map( A => DATA2(6), ZN => n141);
   U129 : INV_X1 port map( A => DATA2(5), ZN => n142);
   U130 : INV_X1 port map( A => DATA2(4), ZN => n143);
   U131 : INV_X1 port map( A => DATA2(3), ZN => n144);
   U132 : INV_X1 port map( A => DATA2(2), ZN => n145);
   U133 : INV_X1 port map( A => DATA2(1), ZN => n146);
   U134 : INV_X1 port map( A => DATA2(0), ZN => n147);
   U135 : INV_X1 port map( A => n36, ZN => n160);
   U136 : NAND3_X1 port map( A1 => n40, A2 => n41, A3 => n42, ZN => OUTALU(0));
   U137 : AOI22_X1 port map( A1 => N79, A2 => n3, B1 => Y_LOGIC_0_port, B2 => 
                           n4, ZN => n42);
   U138 : NAND3_X1 port map( A1 => FUNC(3), A2 => n43, A3 => FUNC(2), ZN => n39
                           );
   U139 : NAND3_X1 port map( A1 => n44, A2 => n45, A3 => FUNC(1), ZN => n38);
   U140 : NAND3_X1 port map( A1 => n43, A2 => n44, A3 => FUNC(3), ZN => n46);
   U141 : NAND3_X1 port map( A1 => n43, A2 => n47, A3 => FUNC(2), ZN => n37);
   U142 : NOR2_X1 port map( A1 => FUNC(1), A2 => FUNC(0), ZN => n43);
   U143 : NAND2_X1 port map( A1 => OUT_SHIFTER_0_port, A2 => n2, ZN => n41);
   U144 : NAND3_X1 port map( A1 => FUNC(2), A2 => n47, A3 => n49, ZN => n48);
   U145 : INV_X1 port map( A => FUNC(3), ZN => n47);
   U146 : NAND3_X1 port map( A1 => FUNC(3), A2 => n44, A3 => n49, ZN => n36);
   U147 : MUX2_X1 port map( A => n50, B => n51, S => FUNC(3), Z => n40);
   U148 : NAND2_X1 port map( A1 => N112, A2 => U2_U2_Z_0, ZN => n51);
   U149 : AOI22_X1 port map( A1 => n52, A2 => N113, B1 => N111, B2 => U2_U2_Z_0
                           , ZN => n50);
   U150 : AND3_X1 port map( A1 => FUNC(2), A2 => n45, A3 => FUNC(1), ZN => 
                           U2_U2_Z_0);
   U151 : AND2_X1 port map( A1 => n44, A2 => n49, ZN => n52);
   U152 : NOR2_X1 port map( A1 => n45, A2 => FUNC(1), ZN => n49);
   U153 : INV_X1 port map( A => FUNC(0), ZN => n45);
   U154 : INV_X1 port map( A => FUNC(2), ZN => n44);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity EXTENDER_NBIT32_IMM_field_lenght16 is

   port( NOT_EXT_IMM : in std_logic_vector (15 downto 0);  SIGNED_IMM : in 
         std_logic;  EXT_IMM : out std_logic_vector (31 downto 0));

end EXTENDER_NBIT32_IMM_field_lenght16;

architecture SYN_BEHAVIOR of EXTENDER_NBIT32_IMM_field_lenght16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal EXT_IMM_31_port : std_logic;

begin
   EXT_IMM <= ( EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, 
      EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, 
      EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, 
      EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, 
      EXT_IMM_31_port, NOT_EXT_IMM(15), NOT_EXT_IMM(14), NOT_EXT_IMM(13), 
      NOT_EXT_IMM(12), NOT_EXT_IMM(11), NOT_EXT_IMM(10), NOT_EXT_IMM(9), 
      NOT_EXT_IMM(8), NOT_EXT_IMM(7), NOT_EXT_IMM(6), NOT_EXT_IMM(5), 
      NOT_EXT_IMM(4), NOT_EXT_IMM(3), NOT_EXT_IMM(2), NOT_EXT_IMM(1), 
      NOT_EXT_IMM(0) );
   
   U2 : AND2_X1 port map( A1 => SIGNED_IMM, A2 => NOT_EXT_IMM(15), ZN => 
                           EXT_IMM_31_port);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REGISTER_FILE_NBIT32_NREG32 is

   port( CLK, RST, EN, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 :
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0));

end REGISTER_FILE_NBIT32_NREG32;

architecture SYN_BEHAVIOR of REGISTER_FILE_NBIT32_NREG32 is

   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component SELECT_OP
      generic( num_inputs, input_width : integer );
      port( DATA : in std_logic_vector( num_inputs* input_width - 1 downto 0 );
            CONTROL : in std_logic_vector( num_inputs - 1 downto 0 ); Z : out 
            std_logic_vector( input_width - 1 downto 0 ) );
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   signal N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, X_Logic1_port, 
      X_Logic0_port, CLK_port, RD1_port, RD2_port, DATAIN_31_port, 
      DATAIN_30_port, DATAIN_29_port, DATAIN_28_port, DATAIN_27_port, 
      DATAIN_26_port, DATAIN_25_port, DATAIN_24_port, DATAIN_23_port, 
      DATAIN_22_port, DATAIN_21_port, DATAIN_20_port, DATAIN_19_port, 
      DATAIN_18_port, DATAIN_17_port, DATAIN_16_port, DATAIN_15_port, 
      DATAIN_14_port, DATAIN_13_port, DATAIN_12_port, DATAIN_11_port, 
      DATAIN_10_port, DATAIN_9_port, DATAIN_8_port, DATAIN_7_port, 
      DATAIN_6_port, DATAIN_5_port, DATAIN_4_port, DATAIN_3_port, DATAIN_2_port
      , DATAIN_1_port, DATAIN_0_port, OUT1_31_port, OUT1_30_port, OUT1_29_port,
      OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, 
      OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, 
      OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, 
      OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, 
      OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, 
      OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port, OUT2_31_port, 
      OUT2_30_port, OUT2_29_port, OUT2_28_port, OUT2_27_port, OUT2_26_port, 
      OUT2_25_port, OUT2_24_port, OUT2_23_port, OUT2_22_port, OUT2_21_port, 
      OUT2_20_port, OUT2_19_port, OUT2_18_port, OUT2_17_port, OUT2_16_port, 
      OUT2_15_port, OUT2_14_port, OUT2_13_port, OUT2_12_port, OUT2_11_port, 
      OUT2_10_port, OUT2_9_port, OUT2_8_port, OUT2_7_port, OUT2_6_port, 
      OUT2_5_port, OUT2_4_port, OUT2_3_port, OUT2_2_port, OUT2_1_port, 
      OUT2_0_port, REGISTERS_0_31_port, REGISTERS_0_30_port, 
      REGISTERS_0_29_port, REGISTERS_0_28_port, REGISTERS_0_27_port, 
      REGISTERS_0_26_port, REGISTERS_0_25_port, REGISTERS_0_24_port, 
      REGISTERS_0_23_port, REGISTERS_0_22_port, REGISTERS_0_21_port, 
      REGISTERS_0_20_port, REGISTERS_0_19_port, REGISTERS_0_18_port, 
      REGISTERS_0_17_port, REGISTERS_0_16_port, REGISTERS_0_15_port, 
      REGISTERS_0_14_port, REGISTERS_0_13_port, REGISTERS_0_12_port, 
      REGISTERS_0_11_port, REGISTERS_0_10_port, REGISTERS_0_9_port, 
      REGISTERS_0_8_port, REGISTERS_0_7_port, REGISTERS_0_6_port, 
      REGISTERS_0_5_port, REGISTERS_0_4_port, REGISTERS_0_3_port, 
      REGISTERS_0_2_port, REGISTERS_0_1_port, REGISTERS_0_0_port, 
      REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_31_port, 
      REGISTERS_2_30_port, REGISTERS_2_29_port, REGISTERS_2_28_port, 
      REGISTERS_2_27_port, REGISTERS_2_26_port, REGISTERS_2_25_port, 
      REGISTERS_2_24_port, REGISTERS_2_23_port, REGISTERS_2_22_port, 
      REGISTERS_2_21_port, REGISTERS_2_20_port, REGISTERS_2_19_port, 
      REGISTERS_2_18_port, REGISTERS_2_17_port, REGISTERS_2_16_port, 
      REGISTERS_2_15_port, REGISTERS_2_14_port, REGISTERS_2_13_port, 
      REGISTERS_2_12_port, REGISTERS_2_11_port, REGISTERS_2_10_port, 
      REGISTERS_2_9_port, REGISTERS_2_8_port, REGISTERS_2_7_port, 
      REGISTERS_2_6_port, REGISTERS_2_5_port, REGISTERS_2_4_port, 
      REGISTERS_2_3_port, REGISTERS_2_2_port, REGISTERS_2_1_port, 
      REGISTERS_2_0_port, REGISTERS_3_31_port, REGISTERS_3_30_port, 
      REGISTERS_3_29_port, REGISTERS_3_28_port, REGISTERS_3_27_port, 
      REGISTERS_3_26_port, REGISTERS_3_25_port, REGISTERS_3_24_port, 
      REGISTERS_3_23_port, REGISTERS_3_22_port, REGISTERS_3_21_port, 
      REGISTERS_3_20_port, REGISTERS_3_19_port, REGISTERS_3_18_port, 
      REGISTERS_3_17_port, REGISTERS_3_16_port, REGISTERS_3_15_port, 
      REGISTERS_3_14_port, REGISTERS_3_13_port, REGISTERS_3_12_port, 
      REGISTERS_3_11_port, REGISTERS_3_10_port, REGISTERS_3_9_port, 
      REGISTERS_3_8_port, REGISTERS_3_7_port, REGISTERS_3_6_port, 
      REGISTERS_3_5_port, REGISTERS_3_4_port, REGISTERS_3_3_port, 
      REGISTERS_3_2_port, REGISTERS_3_1_port, REGISTERS_3_0_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_31_port, 
      REGISTERS_5_30_port, REGISTERS_5_29_port, REGISTERS_5_28_port, 
      REGISTERS_5_27_port, REGISTERS_5_26_port, REGISTERS_5_25_port, 
      REGISTERS_5_24_port, REGISTERS_5_23_port, REGISTERS_5_22_port, 
      REGISTERS_5_21_port, REGISTERS_5_20_port, REGISTERS_5_19_port, 
      REGISTERS_5_18_port, REGISTERS_5_17_port, REGISTERS_5_16_port, 
      REGISTERS_5_15_port, REGISTERS_5_14_port, REGISTERS_5_13_port, 
      REGISTERS_5_12_port, REGISTERS_5_11_port, REGISTERS_5_10_port, 
      REGISTERS_5_9_port, REGISTERS_5_8_port, REGISTERS_5_7_port, 
      REGISTERS_5_6_port, REGISTERS_5_5_port, REGISTERS_5_4_port, 
      REGISTERS_5_3_port, REGISTERS_5_2_port, REGISTERS_5_1_port, 
      REGISTERS_5_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_31_port, 
      REGISTERS_8_30_port, REGISTERS_8_29_port, REGISTERS_8_28_port, 
      REGISTERS_8_27_port, REGISTERS_8_26_port, REGISTERS_8_25_port, 
      REGISTERS_8_24_port, REGISTERS_8_23_port, REGISTERS_8_22_port, 
      REGISTERS_8_21_port, REGISTERS_8_20_port, REGISTERS_8_19_port, 
      REGISTERS_8_18_port, REGISTERS_8_17_port, REGISTERS_8_16_port, 
      REGISTERS_8_15_port, REGISTERS_8_14_port, REGISTERS_8_13_port, 
      REGISTERS_8_12_port, REGISTERS_8_11_port, REGISTERS_8_10_port, 
      REGISTERS_8_9_port, REGISTERS_8_8_port, REGISTERS_8_7_port, 
      REGISTERS_8_6_port, REGISTERS_8_5_port, REGISTERS_8_4_port, 
      REGISTERS_8_3_port, REGISTERS_8_2_port, REGISTERS_8_1_port, 
      REGISTERS_8_0_port, REGISTERS_9_31_port, REGISTERS_9_30_port, 
      REGISTERS_9_29_port, REGISTERS_9_28_port, REGISTERS_9_27_port, 
      REGISTERS_9_26_port, REGISTERS_9_25_port, REGISTERS_9_24_port, 
      REGISTERS_9_23_port, REGISTERS_9_22_port, REGISTERS_9_21_port, 
      REGISTERS_9_20_port, REGISTERS_9_19_port, REGISTERS_9_18_port, 
      REGISTERS_9_17_port, REGISTERS_9_16_port, REGISTERS_9_15_port, 
      REGISTERS_9_14_port, REGISTERS_9_13_port, REGISTERS_9_12_port, 
      REGISTERS_9_11_port, REGISTERS_9_10_port, REGISTERS_9_9_port, 
      REGISTERS_9_8_port, REGISTERS_9_7_port, REGISTERS_9_6_port, 
      REGISTERS_9_5_port, REGISTERS_9_4_port, REGISTERS_9_3_port, 
      REGISTERS_9_2_port, REGISTERS_9_1_port, REGISTERS_9_0_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_31_port, 
      REGISTERS_11_30_port, REGISTERS_11_29_port, REGISTERS_11_28_port, 
      REGISTERS_11_27_port, REGISTERS_11_26_port, REGISTERS_11_25_port, 
      REGISTERS_11_24_port, REGISTERS_11_23_port, REGISTERS_11_22_port, 
      REGISTERS_11_21_port, REGISTERS_11_20_port, REGISTERS_11_19_port, 
      REGISTERS_11_18_port, REGISTERS_11_17_port, REGISTERS_11_16_port, 
      REGISTERS_11_15_port, REGISTERS_11_14_port, REGISTERS_11_13_port, 
      REGISTERS_11_12_port, REGISTERS_11_11_port, REGISTERS_11_10_port, 
      REGISTERS_11_9_port, REGISTERS_11_8_port, REGISTERS_11_7_port, 
      REGISTERS_11_6_port, REGISTERS_11_5_port, REGISTERS_11_4_port, 
      REGISTERS_11_3_port, REGISTERS_11_2_port, REGISTERS_11_1_port, 
      REGISTERS_11_0_port, REGISTERS_12_31_port, REGISTERS_12_30_port, 
      REGISTERS_12_29_port, REGISTERS_12_28_port, REGISTERS_12_27_port, 
      REGISTERS_12_26_port, REGISTERS_12_25_port, REGISTERS_12_24_port, 
      REGISTERS_12_23_port, REGISTERS_12_22_port, REGISTERS_12_21_port, 
      REGISTERS_12_20_port, REGISTERS_12_19_port, REGISTERS_12_18_port, 
      REGISTERS_12_17_port, REGISTERS_12_16_port, REGISTERS_12_15_port, 
      REGISTERS_12_14_port, REGISTERS_12_13_port, REGISTERS_12_12_port, 
      REGISTERS_12_11_port, REGISTERS_12_10_port, REGISTERS_12_9_port, 
      REGISTERS_12_8_port, REGISTERS_12_7_port, REGISTERS_12_6_port, 
      REGISTERS_12_5_port, REGISTERS_12_4_port, REGISTERS_12_3_port, 
      REGISTERS_12_2_port, REGISTERS_12_1_port, REGISTERS_12_0_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_31_port, 
      REGISTERS_14_30_port, REGISTERS_14_29_port, REGISTERS_14_28_port, 
      REGISTERS_14_27_port, REGISTERS_14_26_port, REGISTERS_14_25_port, 
      REGISTERS_14_24_port, REGISTERS_14_23_port, REGISTERS_14_22_port, 
      REGISTERS_14_21_port, REGISTERS_14_20_port, REGISTERS_14_19_port, 
      REGISTERS_14_18_port, REGISTERS_14_17_port, REGISTERS_14_16_port, 
      REGISTERS_14_15_port, REGISTERS_14_14_port, REGISTERS_14_13_port, 
      REGISTERS_14_12_port, REGISTERS_14_11_port, REGISTERS_14_10_port, 
      REGISTERS_14_9_port, REGISTERS_14_8_port, REGISTERS_14_7_port, 
      REGISTERS_14_6_port, REGISTERS_14_5_port, REGISTERS_14_4_port, 
      REGISTERS_14_3_port, REGISTERS_14_2_port, REGISTERS_14_1_port, 
      REGISTERS_14_0_port, REGISTERS_15_31_port, REGISTERS_15_30_port, 
      REGISTERS_15_29_port, REGISTERS_15_28_port, REGISTERS_15_27_port, 
      REGISTERS_15_26_port, REGISTERS_15_25_port, REGISTERS_15_24_port, 
      REGISTERS_15_23_port, REGISTERS_15_22_port, REGISTERS_15_21_port, 
      REGISTERS_15_20_port, REGISTERS_15_19_port, REGISTERS_15_18_port, 
      REGISTERS_15_17_port, REGISTERS_15_16_port, REGISTERS_15_15_port, 
      REGISTERS_15_14_port, REGISTERS_15_13_port, REGISTERS_15_12_port, 
      REGISTERS_15_11_port, REGISTERS_15_10_port, REGISTERS_15_9_port, 
      REGISTERS_15_8_port, REGISTERS_15_7_port, REGISTERS_15_6_port, 
      REGISTERS_15_5_port, REGISTERS_15_4_port, REGISTERS_15_3_port, 
      REGISTERS_15_2_port, REGISTERS_15_1_port, REGISTERS_15_0_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_31_port, 
      REGISTERS_17_30_port, REGISTERS_17_29_port, REGISTERS_17_28_port, 
      REGISTERS_17_27_port, REGISTERS_17_26_port, REGISTERS_17_25_port, 
      REGISTERS_17_24_port, REGISTERS_17_23_port, REGISTERS_17_22_port, 
      REGISTERS_17_21_port, REGISTERS_17_20_port, REGISTERS_17_19_port, 
      REGISTERS_17_18_port, REGISTERS_17_17_port, REGISTERS_17_16_port, 
      REGISTERS_17_15_port, REGISTERS_17_14_port, REGISTERS_17_13_port, 
      REGISTERS_17_12_port, REGISTERS_17_11_port, REGISTERS_17_10_port, 
      REGISTERS_17_9_port, REGISTERS_17_8_port, REGISTERS_17_7_port, 
      REGISTERS_17_6_port, REGISTERS_17_5_port, REGISTERS_17_4_port, 
      REGISTERS_17_3_port, REGISTERS_17_2_port, REGISTERS_17_1_port, 
      REGISTERS_17_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_31_port, 
      REGISTERS_20_30_port, REGISTERS_20_29_port, REGISTERS_20_28_port, 
      REGISTERS_20_27_port, REGISTERS_20_26_port, REGISTERS_20_25_port, 
      REGISTERS_20_24_port, REGISTERS_20_23_port, REGISTERS_20_22_port, 
      REGISTERS_20_21_port, REGISTERS_20_20_port, REGISTERS_20_19_port, 
      REGISTERS_20_18_port, REGISTERS_20_17_port, REGISTERS_20_16_port, 
      REGISTERS_20_15_port, REGISTERS_20_14_port, REGISTERS_20_13_port, 
      REGISTERS_20_12_port, REGISTERS_20_11_port, REGISTERS_20_10_port, 
      REGISTERS_20_9_port, REGISTERS_20_8_port, REGISTERS_20_7_port, 
      REGISTERS_20_6_port, REGISTERS_20_5_port, REGISTERS_20_4_port, 
      REGISTERS_20_3_port, REGISTERS_20_2_port, REGISTERS_20_1_port, 
      REGISTERS_20_0_port, REGISTERS_21_31_port, REGISTERS_21_30_port, 
      REGISTERS_21_29_port, REGISTERS_21_28_port, REGISTERS_21_27_port, 
      REGISTERS_21_26_port, REGISTERS_21_25_port, REGISTERS_21_24_port, 
      REGISTERS_21_23_port, REGISTERS_21_22_port, REGISTERS_21_21_port, 
      REGISTERS_21_20_port, REGISTERS_21_19_port, REGISTERS_21_18_port, 
      REGISTERS_21_17_port, REGISTERS_21_16_port, REGISTERS_21_15_port, 
      REGISTERS_21_14_port, REGISTERS_21_13_port, REGISTERS_21_12_port, 
      REGISTERS_21_11_port, REGISTERS_21_10_port, REGISTERS_21_9_port, 
      REGISTERS_21_8_port, REGISTERS_21_7_port, REGISTERS_21_6_port, 
      REGISTERS_21_5_port, REGISTERS_21_4_port, REGISTERS_21_3_port, 
      REGISTERS_21_2_port, REGISTERS_21_1_port, REGISTERS_21_0_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_31_port, 
      REGISTERS_23_30_port, REGISTERS_23_29_port, REGISTERS_23_28_port, 
      REGISTERS_23_27_port, REGISTERS_23_26_port, REGISTERS_23_25_port, 
      REGISTERS_23_24_port, REGISTERS_23_23_port, REGISTERS_23_22_port, 
      REGISTERS_23_21_port, REGISTERS_23_20_port, REGISTERS_23_19_port, 
      REGISTERS_23_18_port, REGISTERS_23_17_port, REGISTERS_23_16_port, 
      REGISTERS_23_15_port, REGISTERS_23_14_port, REGISTERS_23_13_port, 
      REGISTERS_23_12_port, REGISTERS_23_11_port, REGISTERS_23_10_port, 
      REGISTERS_23_9_port, REGISTERS_23_8_port, REGISTERS_23_7_port, 
      REGISTERS_23_6_port, REGISTERS_23_5_port, REGISTERS_23_4_port, 
      REGISTERS_23_3_port, REGISTERS_23_2_port, REGISTERS_23_1_port, 
      REGISTERS_23_0_port, REGISTERS_24_31_port, REGISTERS_24_30_port, 
      REGISTERS_24_29_port, REGISTERS_24_28_port, REGISTERS_24_27_port, 
      REGISTERS_24_26_port, REGISTERS_24_25_port, REGISTERS_24_24_port, 
      REGISTERS_24_23_port, REGISTERS_24_22_port, REGISTERS_24_21_port, 
      REGISTERS_24_20_port, REGISTERS_24_19_port, REGISTERS_24_18_port, 
      REGISTERS_24_17_port, REGISTERS_24_16_port, REGISTERS_24_15_port, 
      REGISTERS_24_14_port, REGISTERS_24_13_port, REGISTERS_24_12_port, 
      REGISTERS_24_11_port, REGISTERS_24_10_port, REGISTERS_24_9_port, 
      REGISTERS_24_8_port, REGISTERS_24_7_port, REGISTERS_24_6_port, 
      REGISTERS_24_5_port, REGISTERS_24_4_port, REGISTERS_24_3_port, 
      REGISTERS_24_2_port, REGISTERS_24_1_port, REGISTERS_24_0_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_31_port, 
      REGISTERS_26_30_port, REGISTERS_26_29_port, REGISTERS_26_28_port, 
      REGISTERS_26_27_port, REGISTERS_26_26_port, REGISTERS_26_25_port, 
      REGISTERS_26_24_port, REGISTERS_26_23_port, REGISTERS_26_22_port, 
      REGISTERS_26_21_port, REGISTERS_26_20_port, REGISTERS_26_19_port, 
      REGISTERS_26_18_port, REGISTERS_26_17_port, REGISTERS_26_16_port, 
      REGISTERS_26_15_port, REGISTERS_26_14_port, REGISTERS_26_13_port, 
      REGISTERS_26_12_port, REGISTERS_26_11_port, REGISTERS_26_10_port, 
      REGISTERS_26_9_port, REGISTERS_26_8_port, REGISTERS_26_7_port, 
      REGISTERS_26_6_port, REGISTERS_26_5_port, REGISTERS_26_4_port, 
      REGISTERS_26_3_port, REGISTERS_26_2_port, REGISTERS_26_1_port, 
      REGISTERS_26_0_port, REGISTERS_27_31_port, REGISTERS_27_30_port, 
      REGISTERS_27_29_port, REGISTERS_27_28_port, REGISTERS_27_27_port, 
      REGISTERS_27_26_port, REGISTERS_27_25_port, REGISTERS_27_24_port, 
      REGISTERS_27_23_port, REGISTERS_27_22_port, REGISTERS_27_21_port, 
      REGISTERS_27_20_port, REGISTERS_27_19_port, REGISTERS_27_18_port, 
      REGISTERS_27_17_port, REGISTERS_27_16_port, REGISTERS_27_15_port, 
      REGISTERS_27_14_port, REGISTERS_27_13_port, REGISTERS_27_12_port, 
      REGISTERS_27_11_port, REGISTERS_27_10_port, REGISTERS_27_9_port, 
      REGISTERS_27_8_port, REGISTERS_27_7_port, REGISTERS_27_6_port, 
      REGISTERS_27_5_port, REGISTERS_27_4_port, REGISTERS_27_3_port, 
      REGISTERS_27_2_port, REGISTERS_27_1_port, REGISTERS_27_0_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_31_port, 
      REGISTERS_29_30_port, REGISTERS_29_29_port, REGISTERS_29_28_port, 
      REGISTERS_29_27_port, REGISTERS_29_26_port, REGISTERS_29_25_port, 
      REGISTERS_29_24_port, REGISTERS_29_23_port, REGISTERS_29_22_port, 
      REGISTERS_29_21_port, REGISTERS_29_20_port, REGISTERS_29_19_port, 
      REGISTERS_29_18_port, REGISTERS_29_17_port, REGISTERS_29_16_port, 
      REGISTERS_29_15_port, REGISTERS_29_14_port, REGISTERS_29_13_port, 
      REGISTERS_29_12_port, REGISTERS_29_11_port, REGISTERS_29_10_port, 
      REGISTERS_29_9_port, REGISTERS_29_8_port, REGISTERS_29_7_port, 
      REGISTERS_29_6_port, REGISTERS_29_5_port, REGISTERS_29_4_port, 
      REGISTERS_29_3_port, REGISTERS_29_2_port, REGISTERS_29_1_port, 
      REGISTERS_29_0_port, REGISTERS_30_31_port, REGISTERS_30_30_port, 
      REGISTERS_30_29_port, REGISTERS_30_28_port, REGISTERS_30_27_port, 
      REGISTERS_30_26_port, REGISTERS_30_25_port, REGISTERS_30_24_port, 
      REGISTERS_30_23_port, REGISTERS_30_22_port, REGISTERS_30_21_port, 
      REGISTERS_30_20_port, REGISTERS_30_19_port, REGISTERS_30_18_port, 
      REGISTERS_30_17_port, REGISTERS_30_16_port, REGISTERS_30_15_port, 
      REGISTERS_30_14_port, REGISTERS_30_13_port, REGISTERS_30_12_port, 
      REGISTERS_30_11_port, REGISTERS_30_10_port, REGISTERS_30_9_port, 
      REGISTERS_30_8_port, REGISTERS_30_7_port, REGISTERS_30_6_port, 
      REGISTERS_30_5_port, REGISTERS_30_4_port, REGISTERS_30_3_port, 
      REGISTERS_30_2_port, REGISTERS_30_1_port, REGISTERS_30_0_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, N12, N13, N14, N15, N16, N17, 
      N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32
      , N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, 
      N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61
      , N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, 
      N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90
      , N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, 
      N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, 
      N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, 
      N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, 
      N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, 
      N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, 
      N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, 
      N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, 
      N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, 
      N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, 
      N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, 
      N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, 
      N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, 
      N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, 
      N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, 
      N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, 
      N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, 
      N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, 
      N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, 
      N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, 
      N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, 
      N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, 
      N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, 
      N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, 
      N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, 
      N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, 
      N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, 
      N416, N417, N418, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060,
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, 
      n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, 
      n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, 
      n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, 
      n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, 
      n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, 
      n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, 
      n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, 
      n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, 
      n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, 
      n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, 
      n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, 
      n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, 
      n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, 
      n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, 
      n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, 
      n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, 
      n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, 
      n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, 
      n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, 
      n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, 
      n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, 
      n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, 
      n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, 
      n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, 
      n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, 
      n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, 
      n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, 
      n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, 
      n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, 
      n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, 
      n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, 
      n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, 
      n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, 
      n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, 
      n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, 
      n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, 
      n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, 
      n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, 
      n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, 
      n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, 
      n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, 
      n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, 
      n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, 
      n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, 
      n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, 
      n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, 
      n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, 
      n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, 
      n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, 
      n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, 
      n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, 
      n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, 
      n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, 
      n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, 
      n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, 
      n_2141 : std_logic;

begin
   CLK_port <= CLK;
   RD1_port <= RD1;
   RD2_port <= RD2;
   ( DATAIN_31_port, DATAIN_30_port, DATAIN_29_port, DATAIN_28_port, 
      DATAIN_27_port, DATAIN_26_port, DATAIN_25_port, DATAIN_24_port, 
      DATAIN_23_port, DATAIN_22_port, DATAIN_21_port, DATAIN_20_port, 
      DATAIN_19_port, DATAIN_18_port, DATAIN_17_port, DATAIN_16_port, 
      DATAIN_15_port, DATAIN_14_port, DATAIN_13_port, DATAIN_12_port, 
      DATAIN_11_port, DATAIN_10_port, DATAIN_9_port, DATAIN_8_port, 
      DATAIN_7_port, DATAIN_6_port, DATAIN_5_port, DATAIN_4_port, DATAIN_3_port
      , DATAIN_2_port, DATAIN_1_port, DATAIN_0_port ) <= DATAIN;
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   C79_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_31_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_31_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_31_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_31_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_31_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_31_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_31_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_31_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_31_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_31_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_31_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_31_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_31_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_31_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_31_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_31_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_31_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_31_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_31_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_31_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_31_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_31_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_31_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_31_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_31_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_31_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_31_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_31_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_31_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_31_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_31_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_31_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N77 );
   C80_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_30_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_30_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_30_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_30_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_30_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_30_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_30_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_30_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_30_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_30_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_30_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_30_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_30_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_30_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_30_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_30_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_30_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_30_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_30_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_30_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_30_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_30_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_30_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_30_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_30_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_30_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_30_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_30_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_30_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_30_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_30_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_30_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N78 );
   C81_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_29_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_29_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_29_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_29_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_29_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_29_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_29_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_29_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_29_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_29_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_29_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_29_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_29_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_29_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_29_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_29_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_29_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_29_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_29_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_29_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_29_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_29_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_29_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_29_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_29_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_29_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_29_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_29_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_29_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_29_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_29_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_29_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N79 );
   C82_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_28_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_28_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_28_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_28_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_28_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_28_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_28_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_28_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_28_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_28_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_28_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_28_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_28_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_28_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_28_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_28_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_28_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_28_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_28_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_28_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_28_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_28_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_28_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_28_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_28_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_28_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_28_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_28_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_28_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_28_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_28_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_28_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N80 );
   C83_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_27_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_27_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_27_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_27_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_27_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_27_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_27_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_27_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_27_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_27_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_27_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_27_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_27_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_27_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_27_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_27_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_27_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_27_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_27_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_27_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_27_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_27_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_27_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_27_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_27_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_27_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_27_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_27_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_27_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_27_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_27_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_27_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N81 );
   C84_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_26_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_26_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_26_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_26_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_26_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_26_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_26_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_26_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_26_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_26_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_26_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_26_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_26_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_26_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_26_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_26_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_26_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_26_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_26_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_26_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_26_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_26_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_26_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_26_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_26_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_26_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_26_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_26_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_26_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_26_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_26_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_26_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N82 );
   C85_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_25_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_25_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_25_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_25_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_25_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_25_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_25_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_25_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_25_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_25_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_25_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_25_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_25_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_25_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_25_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_25_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_25_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_25_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_25_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_25_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_25_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_25_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_25_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_25_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_25_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_25_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_25_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_25_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_25_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_25_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_25_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_25_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N83 );
   C86_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_24_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_24_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_24_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_24_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_24_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_24_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_24_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_24_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_24_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_24_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_24_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_24_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_24_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_24_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_24_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_24_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_24_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_24_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_24_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_24_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_24_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_24_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_24_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_24_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_24_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_24_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_24_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_24_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_24_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_24_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_24_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_24_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N84 );
   C87_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_23_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_23_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_23_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_23_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_23_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_23_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_23_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_23_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_23_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_23_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_23_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_23_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_23_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_23_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_23_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_23_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_23_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_23_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_23_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_23_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_23_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_23_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_23_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_23_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_23_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_23_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_23_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_23_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_23_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_23_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_23_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_23_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N85 );
   C88_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_22_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_22_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_22_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_22_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_22_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_22_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_22_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_22_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_22_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_22_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_22_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_22_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_22_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_22_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_22_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_22_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_22_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_22_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_22_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_22_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_22_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_22_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_22_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_22_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_22_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_22_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_22_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_22_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_22_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_22_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_22_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_22_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N86 );
   C89_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_21_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_21_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_21_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_21_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_21_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_21_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_21_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_21_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_21_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_21_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_21_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_21_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_21_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_21_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_21_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_21_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_21_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_21_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_21_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_21_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_21_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_21_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_21_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_21_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_21_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_21_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_21_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_21_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_21_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_21_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_21_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_21_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N87 );
   C90_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_20_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_20_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_20_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_20_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_20_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_20_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_20_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_20_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_20_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_20_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_20_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_20_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_20_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_20_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_20_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_20_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_20_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_20_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_20_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_20_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_20_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_20_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_20_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_20_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_20_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_20_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_20_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_20_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_20_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_20_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_20_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_20_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N88 );
   C91_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_19_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_19_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_19_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_19_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_19_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_19_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_19_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_19_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_19_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_19_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_19_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_19_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_19_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_19_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_19_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_19_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_19_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_19_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_19_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_19_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_19_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_19_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_19_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_19_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_19_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_19_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_19_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_19_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_19_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_19_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_19_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_19_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N89 );
   C92_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_18_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_18_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_18_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_18_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_18_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_18_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_18_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_18_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_18_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_18_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_18_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_18_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_18_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_18_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_18_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_18_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_18_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_18_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_18_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_18_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_18_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_18_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_18_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_18_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_18_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_18_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_18_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_18_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_18_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_18_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_18_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_18_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N90 );
   C93_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_17_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_17_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_17_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_17_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_17_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_17_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_17_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_17_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_17_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_17_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_17_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_17_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_17_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_17_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_17_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_17_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_17_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_17_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_17_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_17_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_17_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_17_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_17_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_17_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_17_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_17_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_17_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_17_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_17_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_17_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_17_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_17_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N91 );
   C94_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_16_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_16_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_16_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_16_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_16_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_16_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_16_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_16_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_16_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_16_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_16_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_16_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_16_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_16_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_16_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_16_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_16_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_16_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_16_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_16_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_16_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_16_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_16_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_16_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_16_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_16_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_16_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_16_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_16_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_16_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_16_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_16_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N92 );
   C95_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_15_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_15_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_15_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_15_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_15_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_15_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_15_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_15_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_15_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_15_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_15_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_15_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_15_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_15_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_15_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_15_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_15_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_15_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_15_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_15_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_15_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_15_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_15_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_15_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_15_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_15_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_15_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_15_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_15_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_15_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_15_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_15_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N93 );
   C96_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_14_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_14_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_14_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_14_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_14_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_14_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_14_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_14_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_14_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_14_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_14_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_14_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_14_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_14_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_14_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_14_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_14_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_14_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_14_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_14_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_14_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_14_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_14_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_14_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_14_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_14_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_14_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_14_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_14_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_14_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_14_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_14_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N94 );
   C97_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_13_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_13_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_13_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_13_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_13_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_13_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_13_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_13_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_13_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_13_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_13_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_13_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_13_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_13_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_13_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_13_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_13_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_13_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_13_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_13_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_13_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_13_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_13_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_13_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_13_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_13_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_13_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_13_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_13_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_13_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_13_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_13_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N95 );
   C98_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_12_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_12_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_12_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_12_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_12_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_12_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_12_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_12_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_12_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_12_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_12_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_12_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_12_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_12_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_12_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_12_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_12_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_12_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_12_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_12_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_12_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_12_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_12_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_12_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_12_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_12_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_12_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_12_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_12_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_12_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_12_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_12_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N96 );
   C99_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_11_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_11_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_11_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_11_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_11_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_11_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_11_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_11_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_11_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_11_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_11_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_11_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_11_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_11_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_11_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_11_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_11_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_11_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_11_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_11_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_11_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_11_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_11_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_11_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_11_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_11_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_11_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_11_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_11_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_11_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_11_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_11_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N97 );
   C100_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_10_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_10_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_10_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_10_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_10_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_10_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_10_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_10_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_10_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_10_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_10_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_10_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_10_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_10_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_10_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_10_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_10_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_10_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_10_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_10_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_10_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_10_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_10_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_10_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_10_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_10_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_10_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_10_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_10_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_10_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_10_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_10_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N98 );
   C101_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_9_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_9_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_9_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_9_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_9_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_9_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_9_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_9_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_9_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_9_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_9_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_9_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_9_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_9_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_9_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_9_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_9_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_9_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_9_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_9_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_9_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_9_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_9_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_9_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_9_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_9_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_9_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_9_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_9_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_9_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_9_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_9_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N99 );
   C102_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_8_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_8_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_8_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_8_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_8_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_8_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_8_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_8_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_8_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_8_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_8_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_8_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_8_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_8_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_8_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_8_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_8_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_8_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_8_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_8_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_8_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_8_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_8_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_8_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_8_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_8_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_8_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_8_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_8_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_8_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_8_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_8_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N100 );
   C103_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_7_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_7_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_7_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_7_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_7_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_7_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_7_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_7_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_7_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_7_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_7_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_7_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_7_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_7_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_7_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_7_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_7_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_7_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_7_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_7_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_7_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_7_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_7_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_7_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_7_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_7_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_7_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_7_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_7_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_7_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_7_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_7_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N101 );
   C104_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_6_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_6_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_6_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_6_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_6_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_6_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_6_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_6_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_6_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_6_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_6_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_6_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_6_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_6_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_6_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_6_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_6_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_6_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_6_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_6_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_6_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_6_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_6_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_6_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_6_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_6_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_6_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_6_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_6_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_6_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_6_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_6_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N102 );
   C105_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_5_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_5_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_5_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_5_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_5_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_5_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_5_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_5_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_5_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_5_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_5_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_5_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_5_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_5_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_5_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_5_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_5_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_5_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_5_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_5_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_5_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_5_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_5_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_5_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_5_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_5_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_5_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_5_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_5_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_5_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_5_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_5_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N103 );
   C106_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_4_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_4_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_4_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_4_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_4_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_4_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_4_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_4_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_4_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_4_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_4_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_4_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_4_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_4_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_4_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_4_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_4_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_4_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_4_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_4_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_4_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_4_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_4_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_4_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_4_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_4_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_4_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_4_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_4_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_4_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_4_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_4_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N104 );
   C107_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_3_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_3_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_3_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_3_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_3_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_3_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_3_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_3_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_3_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_3_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_3_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_3_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_3_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_3_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_3_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_3_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_3_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_3_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_3_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_3_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_3_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_3_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_3_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_3_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_3_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_3_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_3_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_3_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_3_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_3_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_3_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_3_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N105 );
   C108_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_2_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_2_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_2_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_2_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_2_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_2_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_2_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_2_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_2_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_2_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_2_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_2_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_2_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_2_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_2_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_2_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_2_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_2_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_2_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_2_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_2_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_2_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_2_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_2_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_2_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_2_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_2_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_2_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_2_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_2_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_2_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_2_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N106 );
   C109_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_1_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_1_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_1_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_1_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_1_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_1_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_1_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_1_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_1_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_1_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_1_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_1_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_1_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_1_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_1_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_1_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_1_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_1_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_1_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_1_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_1_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_1_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N107 );
   C110_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_0_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_0_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_0_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_0_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_0_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_0_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_0_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_0_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_0_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_0_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_0_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_0_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_0_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_0_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_0_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_0_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N49, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N53, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N55, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N57, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N59, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N61, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N63, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N65, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N67, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N69, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N71, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N73, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N75, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N46, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N48, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N50, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N52, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N54, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N56, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N58, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N60, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N62, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N64, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N66, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N68, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N70, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N72, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N74, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N76, 
         -- Connections to port 'Z'
         Z(0) => N108 );
   C256_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_31_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_31_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_31_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_31_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_31_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_31_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_31_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_31_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_31_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_31_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_31_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_31_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_31_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_31_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_31_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_31_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_31_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_31_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_31_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_31_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_31_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_31_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_31_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_31_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_31_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_31_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_31_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_31_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_31_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_31_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_31_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_31_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N174 );
   C257_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_30_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_30_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_30_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_30_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_30_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_30_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_30_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_30_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_30_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_30_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_30_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_30_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_30_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_30_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_30_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_30_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_30_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_30_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_30_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_30_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_30_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_30_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_30_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_30_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_30_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_30_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_30_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_30_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_30_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_30_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_30_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_30_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N175 );
   C258_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_29_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_29_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_29_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_29_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_29_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_29_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_29_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_29_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_29_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_29_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_29_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_29_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_29_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_29_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_29_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_29_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_29_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_29_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_29_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_29_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_29_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_29_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_29_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_29_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_29_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_29_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_29_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_29_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_29_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_29_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_29_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_29_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N176 );
   C259_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_28_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_28_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_28_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_28_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_28_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_28_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_28_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_28_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_28_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_28_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_28_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_28_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_28_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_28_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_28_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_28_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_28_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_28_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_28_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_28_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_28_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_28_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_28_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_28_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_28_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_28_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_28_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_28_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_28_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_28_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_28_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_28_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N177 );
   C260_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_27_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_27_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_27_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_27_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_27_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_27_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_27_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_27_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_27_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_27_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_27_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_27_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_27_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_27_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_27_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_27_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_27_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_27_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_27_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_27_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_27_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_27_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_27_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_27_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_27_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_27_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_27_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_27_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_27_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_27_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_27_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_27_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N178 );
   C261_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_26_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_26_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_26_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_26_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_26_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_26_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_26_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_26_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_26_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_26_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_26_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_26_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_26_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_26_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_26_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_26_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_26_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_26_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_26_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_26_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_26_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_26_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_26_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_26_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_26_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_26_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_26_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_26_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_26_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_26_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_26_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_26_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N179 );
   C262_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_25_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_25_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_25_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_25_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_25_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_25_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_25_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_25_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_25_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_25_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_25_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_25_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_25_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_25_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_25_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_25_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_25_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_25_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_25_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_25_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_25_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_25_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_25_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_25_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_25_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_25_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_25_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_25_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_25_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_25_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_25_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_25_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N180 );
   C263_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_24_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_24_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_24_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_24_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_24_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_24_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_24_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_24_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_24_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_24_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_24_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_24_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_24_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_24_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_24_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_24_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_24_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_24_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_24_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_24_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_24_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_24_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_24_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_24_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_24_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_24_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_24_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_24_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_24_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_24_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_24_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_24_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N181 );
   C264_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_23_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_23_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_23_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_23_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_23_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_23_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_23_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_23_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_23_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_23_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_23_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_23_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_23_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_23_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_23_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_23_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_23_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_23_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_23_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_23_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_23_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_23_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_23_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_23_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_23_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_23_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_23_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_23_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_23_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_23_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_23_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_23_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N182 );
   C265_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_22_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_22_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_22_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_22_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_22_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_22_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_22_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_22_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_22_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_22_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_22_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_22_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_22_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_22_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_22_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_22_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_22_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_22_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_22_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_22_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_22_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_22_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_22_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_22_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_22_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_22_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_22_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_22_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_22_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_22_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_22_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_22_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N183 );
   C266_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_21_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_21_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_21_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_21_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_21_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_21_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_21_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_21_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_21_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_21_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_21_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_21_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_21_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_21_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_21_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_21_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_21_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_21_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_21_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_21_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_21_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_21_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_21_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_21_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_21_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_21_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_21_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_21_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_21_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_21_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_21_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_21_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N184 );
   C267_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_20_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_20_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_20_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_20_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_20_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_20_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_20_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_20_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_20_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_20_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_20_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_20_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_20_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_20_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_20_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_20_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_20_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_20_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_20_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_20_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_20_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_20_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_20_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_20_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_20_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_20_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_20_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_20_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_20_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_20_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_20_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_20_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N185 );
   C268_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_19_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_19_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_19_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_19_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_19_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_19_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_19_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_19_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_19_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_19_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_19_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_19_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_19_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_19_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_19_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_19_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_19_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_19_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_19_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_19_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_19_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_19_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_19_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_19_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_19_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_19_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_19_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_19_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_19_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_19_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_19_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_19_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N186 );
   C269_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_18_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_18_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_18_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_18_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_18_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_18_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_18_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_18_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_18_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_18_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_18_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_18_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_18_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_18_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_18_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_18_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_18_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_18_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_18_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_18_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_18_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_18_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_18_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_18_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_18_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_18_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_18_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_18_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_18_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_18_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_18_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_18_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N187 );
   C270_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_17_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_17_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_17_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_17_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_17_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_17_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_17_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_17_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_17_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_17_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_17_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_17_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_17_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_17_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_17_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_17_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_17_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_17_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_17_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_17_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_17_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_17_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_17_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_17_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_17_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_17_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_17_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_17_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_17_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_17_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_17_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_17_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N188 );
   C271_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_16_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_16_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_16_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_16_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_16_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_16_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_16_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_16_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_16_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_16_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_16_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_16_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_16_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_16_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_16_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_16_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_16_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_16_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_16_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_16_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_16_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_16_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_16_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_16_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_16_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_16_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_16_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_16_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_16_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_16_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_16_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_16_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N189 );
   C272_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_15_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_15_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_15_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_15_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_15_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_15_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_15_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_15_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_15_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_15_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_15_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_15_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_15_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_15_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_15_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_15_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_15_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_15_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_15_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_15_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_15_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_15_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_15_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_15_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_15_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_15_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_15_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_15_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_15_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_15_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_15_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_15_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N190 );
   C273_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_14_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_14_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_14_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_14_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_14_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_14_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_14_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_14_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_14_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_14_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_14_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_14_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_14_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_14_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_14_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_14_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_14_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_14_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_14_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_14_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_14_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_14_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_14_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_14_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_14_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_14_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_14_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_14_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_14_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_14_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_14_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_14_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N191 );
   C274_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_13_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_13_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_13_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_13_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_13_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_13_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_13_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_13_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_13_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_13_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_13_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_13_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_13_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_13_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_13_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_13_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_13_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_13_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_13_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_13_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_13_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_13_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_13_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_13_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_13_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_13_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_13_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_13_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_13_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_13_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_13_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_13_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N192 );
   C275_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_12_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_12_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_12_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_12_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_12_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_12_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_12_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_12_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_12_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_12_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_12_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_12_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_12_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_12_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_12_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_12_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_12_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_12_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_12_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_12_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_12_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_12_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_12_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_12_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_12_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_12_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_12_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_12_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_12_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_12_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_12_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_12_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N193 );
   C276_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_11_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_11_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_11_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_11_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_11_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_11_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_11_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_11_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_11_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_11_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_11_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_11_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_11_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_11_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_11_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_11_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_11_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_11_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_11_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_11_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_11_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_11_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_11_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_11_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_11_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_11_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_11_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_11_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_11_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_11_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_11_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_11_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N194 );
   C277_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_10_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_10_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_10_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_10_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_10_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_10_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_10_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_10_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_10_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_10_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_10_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_10_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_10_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_10_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_10_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_10_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_10_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_10_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_10_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_10_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_10_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_10_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_10_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_10_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_10_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_10_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_10_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_10_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_10_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_10_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_10_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_10_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N195 );
   C278_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_9_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_9_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_9_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_9_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_9_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_9_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_9_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_9_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_9_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_9_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_9_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_9_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_9_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_9_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_9_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_9_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_9_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_9_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_9_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_9_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_9_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_9_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_9_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_9_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_9_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_9_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_9_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_9_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_9_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_9_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_9_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_9_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N196 );
   C279_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_8_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_8_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_8_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_8_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_8_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_8_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_8_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_8_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_8_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_8_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_8_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_8_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_8_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_8_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_8_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_8_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_8_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_8_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_8_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_8_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_8_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_8_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_8_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_8_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_8_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_8_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_8_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_8_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_8_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_8_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_8_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_8_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N197 );
   C280_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_7_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_7_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_7_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_7_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_7_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_7_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_7_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_7_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_7_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_7_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_7_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_7_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_7_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_7_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_7_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_7_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_7_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_7_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_7_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_7_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_7_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_7_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_7_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_7_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_7_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_7_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_7_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_7_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_7_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_7_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_7_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_7_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N198 );
   C281_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_6_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_6_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_6_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_6_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_6_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_6_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_6_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_6_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_6_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_6_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_6_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_6_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_6_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_6_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_6_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_6_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_6_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_6_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_6_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_6_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_6_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_6_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_6_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_6_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_6_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_6_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_6_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_6_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_6_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_6_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_6_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_6_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N199 );
   C282_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_5_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_5_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_5_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_5_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_5_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_5_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_5_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_5_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_5_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_5_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_5_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_5_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_5_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_5_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_5_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_5_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_5_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_5_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_5_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_5_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_5_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_5_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_5_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_5_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_5_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_5_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_5_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_5_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_5_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_5_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_5_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_5_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N200 );
   C283_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_4_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_4_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_4_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_4_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_4_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_4_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_4_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_4_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_4_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_4_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_4_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_4_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_4_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_4_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_4_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_4_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_4_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_4_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_4_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_4_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_4_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_4_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_4_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_4_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_4_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_4_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_4_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_4_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_4_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_4_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_4_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_4_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N201 );
   C284_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_3_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_3_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_3_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_3_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_3_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_3_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_3_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_3_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_3_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_3_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_3_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_3_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_3_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_3_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_3_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_3_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_3_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_3_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_3_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_3_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_3_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_3_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_3_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_3_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_3_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_3_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_3_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_3_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_3_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_3_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_3_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_3_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N202 );
   C285_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_2_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_2_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_2_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_2_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_2_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_2_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_2_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_2_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_2_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_2_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_2_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_2_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_2_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_2_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_2_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_2_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_2_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_2_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_2_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_2_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_2_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_2_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_2_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_2_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_2_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_2_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_2_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_2_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_2_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_2_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_2_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_2_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N203 );
   C286_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_1_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_1_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_1_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_1_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_1_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_1_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_1_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_1_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_1_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_1_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_1_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_1_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_1_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_1_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_1_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_1_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_1_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_1_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_1_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_1_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_1_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_1_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N204 );
   C287_cell : SELECT_OP
      generic map ( num_inputs => 32, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => REGISTERS_0_0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => REGISTERS_1_0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => REGISTERS_2_0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => REGISTERS_3_0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => REGISTERS_4_0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => REGISTERS_5_0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => REGISTERS_6_0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => REGISTERS_7_0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => REGISTERS_8_0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => REGISTERS_9_0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => REGISTERS_10_0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => REGISTERS_11_0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => REGISTERS_12_0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => REGISTERS_13_0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => REGISTERS_14_0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => REGISTERS_15_0_port, 
         -- Connections to port 'DATA17'
         DATA(16) => REGISTERS_16_0_port, 
         -- Connections to port 'DATA18'
         DATA(17) => REGISTERS_17_0_port, 
         -- Connections to port 'DATA19'
         DATA(18) => REGISTERS_18_0_port, 
         -- Connections to port 'DATA20'
         DATA(19) => REGISTERS_19_0_port, 
         -- Connections to port 'DATA21'
         DATA(20) => REGISTERS_20_0_port, 
         -- Connections to port 'DATA22'
         DATA(21) => REGISTERS_21_0_port, 
         -- Connections to port 'DATA23'
         DATA(22) => REGISTERS_22_0_port, 
         -- Connections to port 'DATA24'
         DATA(23) => REGISTERS_23_0_port, 
         -- Connections to port 'DATA25'
         DATA(24) => REGISTERS_24_0_port, 
         -- Connections to port 'DATA26'
         DATA(25) => REGISTERS_25_0_port, 
         -- Connections to port 'DATA27'
         DATA(26) => REGISTERS_26_0_port, 
         -- Connections to port 'DATA28'
         DATA(27) => REGISTERS_27_0_port, 
         -- Connections to port 'DATA29'
         DATA(28) => REGISTERS_28_0_port, 
         -- Connections to port 'DATA30'
         DATA(29) => REGISTERS_29_0_port, 
         -- Connections to port 'DATA31'
         DATA(30) => REGISTERS_30_0_port, 
         -- Connections to port 'DATA32'
         DATA(31) => REGISTERS_31_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N142, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N144, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N146, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N148, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N150, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N152, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N154, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N156, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N158, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N160, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N162, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N164, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N166, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N168, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N170, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N172, 
         -- Connections to port 'CONTROL17'
         CONTROL(16) => N143, 
         -- Connections to port 'CONTROL18'
         CONTROL(17) => N145, 
         -- Connections to port 'CONTROL19'
         CONTROL(18) => N147, 
         -- Connections to port 'CONTROL20'
         CONTROL(19) => N149, 
         -- Connections to port 'CONTROL21'
         CONTROL(20) => N151, 
         -- Connections to port 'CONTROL22'
         CONTROL(21) => N153, 
         -- Connections to port 'CONTROL23'
         CONTROL(22) => N155, 
         -- Connections to port 'CONTROL24'
         CONTROL(23) => N157, 
         -- Connections to port 'CONTROL25'
         CONTROL(24) => N159, 
         -- Connections to port 'CONTROL26'
         CONTROL(25) => N161, 
         -- Connections to port 'CONTROL27'
         CONTROL(26) => N163, 
         -- Connections to port 'CONTROL28'
         CONTROL(27) => N165, 
         -- Connections to port 'CONTROL29'
         CONTROL(28) => N167, 
         -- Connections to port 'CONTROL30'
         CONTROL(29) => N169, 
         -- Connections to port 'CONTROL31'
         CONTROL(30) => N171, 
         -- Connections to port 'CONTROL32'
         CONTROL(31) => N173, 
         -- Connections to port 'Z'
         Z(0) => N205 );
   REGISTERS_reg_0_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_0_31_port, QN => n_1054);
   REGISTERS_reg_0_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_0_30_port, QN => n_1055);
   REGISTERS_reg_0_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_0_29_port, QN => n_1056);
   REGISTERS_reg_0_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_0_28_port, QN => n_1057);
   REGISTERS_reg_0_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_0_27_port, QN => n_1058);
   REGISTERS_reg_0_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_0_26_port, QN => n_1059);
   REGISTERS_reg_0_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_0_25_port, QN => n_1060);
   REGISTERS_reg_0_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_0_24_port, QN => n_1061);
   REGISTERS_reg_0_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_0_23_port, QN => n_1062);
   REGISTERS_reg_0_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_0_22_port, QN => n_1063);
   REGISTERS_reg_0_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_0_21_port, QN => n_1064);
   REGISTERS_reg_0_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_0_20_port, QN => n_1065);
   REGISTERS_reg_0_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_0_19_port, QN => n_1066);
   REGISTERS_reg_0_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_0_18_port, QN => n_1067);
   REGISTERS_reg_0_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_0_17_port, QN => n_1068);
   REGISTERS_reg_0_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_0_16_port, QN => n_1069);
   REGISTERS_reg_0_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_0_15_port, QN => n_1070);
   REGISTERS_reg_0_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_0_14_port, QN => n_1071);
   REGISTERS_reg_0_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_0_13_port, QN => n_1072);
   REGISTERS_reg_0_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_0_12_port, QN => n_1073);
   REGISTERS_reg_0_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_0_11_port, QN => n_1074);
   REGISTERS_reg_0_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_0_10_port, QN => n_1075);
   REGISTERS_reg_0_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_0_9_port, QN => n_1076);
   REGISTERS_reg_0_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_0_8_port, QN => n_1077);
   REGISTERS_reg_0_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_0_7_port, QN => n_1078);
   REGISTERS_reg_0_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_0_6_port, QN => n_1079);
   REGISTERS_reg_0_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_0_5_port, QN => n_1080);
   REGISTERS_reg_0_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_0_4_port, QN => n_1081);
   REGISTERS_reg_0_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_0_3_port, QN => n_1082);
   REGISTERS_reg_0_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_0_2_port, QN => n_1083);
   REGISTERS_reg_0_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_0_1_port, QN => n_1084);
   REGISTERS_reg_0_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N302, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_0_0_port, QN => n_1085);
   REGISTERS_reg_1_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_1_31_port, QN => n_1086);
   REGISTERS_reg_1_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_1_30_port, QN => n_1087);
   REGISTERS_reg_1_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_1_29_port, QN => n_1088);
   REGISTERS_reg_1_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_1_28_port, QN => n_1089);
   REGISTERS_reg_1_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_1_27_port, QN => n_1090);
   REGISTERS_reg_1_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_1_26_port, QN => n_1091);
   REGISTERS_reg_1_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_1_25_port, QN => n_1092);
   REGISTERS_reg_1_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_1_24_port, QN => n_1093);
   REGISTERS_reg_1_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_1_23_port, QN => n_1094);
   REGISTERS_reg_1_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_1_22_port, QN => n_1095);
   REGISTERS_reg_1_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_1_21_port, QN => n_1096);
   REGISTERS_reg_1_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_1_20_port, QN => n_1097);
   REGISTERS_reg_1_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_1_19_port, QN => n_1098);
   REGISTERS_reg_1_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_1_18_port, QN => n_1099);
   REGISTERS_reg_1_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_1_17_port, QN => n_1100);
   REGISTERS_reg_1_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_1_16_port, QN => n_1101);
   REGISTERS_reg_1_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_1_15_port, QN => n_1102);
   REGISTERS_reg_1_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_1_14_port, QN => n_1103);
   REGISTERS_reg_1_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_1_13_port, QN => n_1104);
   REGISTERS_reg_1_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_1_12_port, QN => n_1105);
   REGISTERS_reg_1_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_1_11_port, QN => n_1106);
   REGISTERS_reg_1_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_1_10_port, QN => n_1107);
   REGISTERS_reg_1_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_1_9_port, QN => n_1108);
   REGISTERS_reg_1_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_1_8_port, QN => n_1109);
   REGISTERS_reg_1_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_1_7_port, QN => n_1110);
   REGISTERS_reg_1_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_1_6_port, QN => n_1111);
   REGISTERS_reg_1_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_1_5_port, QN => n_1112);
   REGISTERS_reg_1_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_1_4_port, QN => n_1113);
   REGISTERS_reg_1_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_1_3_port, QN => n_1114);
   REGISTERS_reg_1_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_1_2_port, QN => n_1115);
   REGISTERS_reg_1_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_1_1_port, QN => n_1116);
   REGISTERS_reg_1_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N301, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_1_0_port, QN => n_1117);
   REGISTERS_reg_2_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_2_31_port, QN => n_1118);
   REGISTERS_reg_2_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_2_30_port, QN => n_1119);
   REGISTERS_reg_2_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_2_29_port, QN => n_1120);
   REGISTERS_reg_2_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_2_28_port, QN => n_1121);
   REGISTERS_reg_2_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_2_27_port, QN => n_1122);
   REGISTERS_reg_2_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_2_26_port, QN => n_1123);
   REGISTERS_reg_2_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_2_25_port, QN => n_1124);
   REGISTERS_reg_2_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_2_24_port, QN => n_1125);
   REGISTERS_reg_2_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_2_23_port, QN => n_1126);
   REGISTERS_reg_2_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_2_22_port, QN => n_1127);
   REGISTERS_reg_2_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_2_21_port, QN => n_1128);
   REGISTERS_reg_2_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_2_20_port, QN => n_1129);
   REGISTERS_reg_2_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_2_19_port, QN => n_1130);
   REGISTERS_reg_2_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_2_18_port, QN => n_1131);
   REGISTERS_reg_2_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_2_17_port, QN => n_1132);
   REGISTERS_reg_2_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_2_16_port, QN => n_1133);
   REGISTERS_reg_2_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_2_15_port, QN => n_1134);
   REGISTERS_reg_2_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_2_14_port, QN => n_1135);
   REGISTERS_reg_2_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_2_13_port, QN => n_1136);
   REGISTERS_reg_2_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_2_12_port, QN => n_1137);
   REGISTERS_reg_2_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_2_11_port, QN => n_1138);
   REGISTERS_reg_2_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_2_10_port, QN => n_1139);
   REGISTERS_reg_2_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_2_9_port, QN => n_1140);
   REGISTERS_reg_2_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_2_8_port, QN => n_1141);
   REGISTERS_reg_2_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_2_7_port, QN => n_1142);
   REGISTERS_reg_2_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_2_6_port, QN => n_1143);
   REGISTERS_reg_2_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_2_5_port, QN => n_1144);
   REGISTERS_reg_2_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_2_4_port, QN => n_1145);
   REGISTERS_reg_2_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_2_3_port, QN => n_1146);
   REGISTERS_reg_2_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_2_2_port, QN => n_1147);
   REGISTERS_reg_2_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_2_1_port, QN => n_1148);
   REGISTERS_reg_2_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N300, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_2_0_port, QN => n_1149);
   REGISTERS_reg_3_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_3_31_port, QN => n_1150);
   REGISTERS_reg_3_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_3_30_port, QN => n_1151);
   REGISTERS_reg_3_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_3_29_port, QN => n_1152);
   REGISTERS_reg_3_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_3_28_port, QN => n_1153);
   REGISTERS_reg_3_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_3_27_port, QN => n_1154);
   REGISTERS_reg_3_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_3_26_port, QN => n_1155);
   REGISTERS_reg_3_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_3_25_port, QN => n_1156);
   REGISTERS_reg_3_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_3_24_port, QN => n_1157);
   REGISTERS_reg_3_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_3_23_port, QN => n_1158);
   REGISTERS_reg_3_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_3_22_port, QN => n_1159);
   REGISTERS_reg_3_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_3_21_port, QN => n_1160);
   REGISTERS_reg_3_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_3_20_port, QN => n_1161);
   REGISTERS_reg_3_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_3_19_port, QN => n_1162);
   REGISTERS_reg_3_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_3_18_port, QN => n_1163);
   REGISTERS_reg_3_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_3_17_port, QN => n_1164);
   REGISTERS_reg_3_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_3_16_port, QN => n_1165);
   REGISTERS_reg_3_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_3_15_port, QN => n_1166);
   REGISTERS_reg_3_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_3_14_port, QN => n_1167);
   REGISTERS_reg_3_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_3_13_port, QN => n_1168);
   REGISTERS_reg_3_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_3_12_port, QN => n_1169);
   REGISTERS_reg_3_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_3_11_port, QN => n_1170);
   REGISTERS_reg_3_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_3_10_port, QN => n_1171);
   REGISTERS_reg_3_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_3_9_port, QN => n_1172);
   REGISTERS_reg_3_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_3_8_port, QN => n_1173);
   REGISTERS_reg_3_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_3_7_port, QN => n_1174);
   REGISTERS_reg_3_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_3_6_port, QN => n_1175);
   REGISTERS_reg_3_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_3_5_port, QN => n_1176);
   REGISTERS_reg_3_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_3_4_port, QN => n_1177);
   REGISTERS_reg_3_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_3_3_port, QN => n_1178);
   REGISTERS_reg_3_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_3_2_port, QN => n_1179);
   REGISTERS_reg_3_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_3_1_port, QN => n_1180);
   REGISTERS_reg_3_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N299, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_3_0_port, QN => n_1181);
   REGISTERS_reg_4_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_4_31_port, QN => n_1182);
   REGISTERS_reg_4_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_4_30_port, QN => n_1183);
   REGISTERS_reg_4_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_4_29_port, QN => n_1184);
   REGISTERS_reg_4_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_4_28_port, QN => n_1185);
   REGISTERS_reg_4_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_4_27_port, QN => n_1186);
   REGISTERS_reg_4_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_4_26_port, QN => n_1187);
   REGISTERS_reg_4_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_4_25_port, QN => n_1188);
   REGISTERS_reg_4_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_4_24_port, QN => n_1189);
   REGISTERS_reg_4_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_4_23_port, QN => n_1190);
   REGISTERS_reg_4_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_4_22_port, QN => n_1191);
   REGISTERS_reg_4_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_4_21_port, QN => n_1192);
   REGISTERS_reg_4_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_4_20_port, QN => n_1193);
   REGISTERS_reg_4_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_4_19_port, QN => n_1194);
   REGISTERS_reg_4_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_4_18_port, QN => n_1195);
   REGISTERS_reg_4_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_4_17_port, QN => n_1196);
   REGISTERS_reg_4_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_4_16_port, QN => n_1197);
   REGISTERS_reg_4_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_4_15_port, QN => n_1198);
   REGISTERS_reg_4_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_4_14_port, QN => n_1199);
   REGISTERS_reg_4_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_4_13_port, QN => n_1200);
   REGISTERS_reg_4_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_4_12_port, QN => n_1201);
   REGISTERS_reg_4_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_4_11_port, QN => n_1202);
   REGISTERS_reg_4_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_4_10_port, QN => n_1203);
   REGISTERS_reg_4_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_4_9_port, QN => n_1204);
   REGISTERS_reg_4_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_4_8_port, QN => n_1205);
   REGISTERS_reg_4_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_4_7_port, QN => n_1206);
   REGISTERS_reg_4_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_4_6_port, QN => n_1207);
   REGISTERS_reg_4_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_4_5_port, QN => n_1208);
   REGISTERS_reg_4_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_4_4_port, QN => n_1209);
   REGISTERS_reg_4_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_4_3_port, QN => n_1210);
   REGISTERS_reg_4_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_4_2_port, QN => n_1211);
   REGISTERS_reg_4_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_4_1_port, QN => n_1212);
   REGISTERS_reg_4_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N298, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_4_0_port, QN => n_1213);
   REGISTERS_reg_5_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_5_31_port, QN => n_1214);
   REGISTERS_reg_5_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_5_30_port, QN => n_1215);
   REGISTERS_reg_5_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_5_29_port, QN => n_1216);
   REGISTERS_reg_5_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_5_28_port, QN => n_1217);
   REGISTERS_reg_5_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_5_27_port, QN => n_1218);
   REGISTERS_reg_5_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_5_26_port, QN => n_1219);
   REGISTERS_reg_5_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_5_25_port, QN => n_1220);
   REGISTERS_reg_5_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_5_24_port, QN => n_1221);
   REGISTERS_reg_5_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_5_23_port, QN => n_1222);
   REGISTERS_reg_5_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_5_22_port, QN => n_1223);
   REGISTERS_reg_5_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_5_21_port, QN => n_1224);
   REGISTERS_reg_5_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_5_20_port, QN => n_1225);
   REGISTERS_reg_5_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_5_19_port, QN => n_1226);
   REGISTERS_reg_5_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_5_18_port, QN => n_1227);
   REGISTERS_reg_5_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_5_17_port, QN => n_1228);
   REGISTERS_reg_5_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_5_16_port, QN => n_1229);
   REGISTERS_reg_5_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_5_15_port, QN => n_1230);
   REGISTERS_reg_5_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_5_14_port, QN => n_1231);
   REGISTERS_reg_5_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_5_13_port, QN => n_1232);
   REGISTERS_reg_5_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_5_12_port, QN => n_1233);
   REGISTERS_reg_5_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_5_11_port, QN => n_1234);
   REGISTERS_reg_5_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_5_10_port, QN => n_1235);
   REGISTERS_reg_5_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_5_9_port, QN => n_1236);
   REGISTERS_reg_5_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_5_8_port, QN => n_1237);
   REGISTERS_reg_5_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_5_7_port, QN => n_1238);
   REGISTERS_reg_5_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_5_6_port, QN => n_1239);
   REGISTERS_reg_5_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_5_5_port, QN => n_1240);
   REGISTERS_reg_5_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_5_4_port, QN => n_1241);
   REGISTERS_reg_5_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_5_3_port, QN => n_1242);
   REGISTERS_reg_5_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_5_2_port, QN => n_1243);
   REGISTERS_reg_5_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_5_1_port, QN => n_1244);
   REGISTERS_reg_5_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N297, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_5_0_port, QN => n_1245);
   REGISTERS_reg_6_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_6_31_port, QN => n_1246);
   REGISTERS_reg_6_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_6_30_port, QN => n_1247);
   REGISTERS_reg_6_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_6_29_port, QN => n_1248);
   REGISTERS_reg_6_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_6_28_port, QN => n_1249);
   REGISTERS_reg_6_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_6_27_port, QN => n_1250);
   REGISTERS_reg_6_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_6_26_port, QN => n_1251);
   REGISTERS_reg_6_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_6_25_port, QN => n_1252);
   REGISTERS_reg_6_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_6_24_port, QN => n_1253);
   REGISTERS_reg_6_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_6_23_port, QN => n_1254);
   REGISTERS_reg_6_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_6_22_port, QN => n_1255);
   REGISTERS_reg_6_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_6_21_port, QN => n_1256);
   REGISTERS_reg_6_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_6_20_port, QN => n_1257);
   REGISTERS_reg_6_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_6_19_port, QN => n_1258);
   REGISTERS_reg_6_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_6_18_port, QN => n_1259);
   REGISTERS_reg_6_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_6_17_port, QN => n_1260);
   REGISTERS_reg_6_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_6_16_port, QN => n_1261);
   REGISTERS_reg_6_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_6_15_port, QN => n_1262);
   REGISTERS_reg_6_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_6_14_port, QN => n_1263);
   REGISTERS_reg_6_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_6_13_port, QN => n_1264);
   REGISTERS_reg_6_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_6_12_port, QN => n_1265);
   REGISTERS_reg_6_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_6_11_port, QN => n_1266);
   REGISTERS_reg_6_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_6_10_port, QN => n_1267);
   REGISTERS_reg_6_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_6_9_port, QN => n_1268);
   REGISTERS_reg_6_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_6_8_port, QN => n_1269);
   REGISTERS_reg_6_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_6_7_port, QN => n_1270);
   REGISTERS_reg_6_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_6_6_port, QN => n_1271);
   REGISTERS_reg_6_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_6_5_port, QN => n_1272);
   REGISTERS_reg_6_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_6_4_port, QN => n_1273);
   REGISTERS_reg_6_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_6_3_port, QN => n_1274);
   REGISTERS_reg_6_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_6_2_port, QN => n_1275);
   REGISTERS_reg_6_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_6_1_port, QN => n_1276);
   REGISTERS_reg_6_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N296, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_6_0_port, QN => n_1277);
   REGISTERS_reg_7_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_7_31_port, QN => n_1278);
   REGISTERS_reg_7_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_7_30_port, QN => n_1279);
   REGISTERS_reg_7_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_7_29_port, QN => n_1280);
   REGISTERS_reg_7_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_7_28_port, QN => n_1281);
   REGISTERS_reg_7_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_7_27_port, QN => n_1282);
   REGISTERS_reg_7_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_7_26_port, QN => n_1283);
   REGISTERS_reg_7_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_7_25_port, QN => n_1284);
   REGISTERS_reg_7_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_7_24_port, QN => n_1285);
   REGISTERS_reg_7_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_7_23_port, QN => n_1286);
   REGISTERS_reg_7_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_7_22_port, QN => n_1287);
   REGISTERS_reg_7_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_7_21_port, QN => n_1288);
   REGISTERS_reg_7_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_7_20_port, QN => n_1289);
   REGISTERS_reg_7_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_7_19_port, QN => n_1290);
   REGISTERS_reg_7_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_7_18_port, QN => n_1291);
   REGISTERS_reg_7_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_7_17_port, QN => n_1292);
   REGISTERS_reg_7_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_7_16_port, QN => n_1293);
   REGISTERS_reg_7_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_7_15_port, QN => n_1294);
   REGISTERS_reg_7_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_7_14_port, QN => n_1295);
   REGISTERS_reg_7_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_7_13_port, QN => n_1296);
   REGISTERS_reg_7_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_7_12_port, QN => n_1297);
   REGISTERS_reg_7_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_7_11_port, QN => n_1298);
   REGISTERS_reg_7_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_7_10_port, QN => n_1299);
   REGISTERS_reg_7_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_7_9_port, QN => n_1300);
   REGISTERS_reg_7_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_7_8_port, QN => n_1301);
   REGISTERS_reg_7_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_7_7_port, QN => n_1302);
   REGISTERS_reg_7_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_7_6_port, QN => n_1303);
   REGISTERS_reg_7_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_7_5_port, QN => n_1304);
   REGISTERS_reg_7_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_7_4_port, QN => n_1305);
   REGISTERS_reg_7_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_7_3_port, QN => n_1306);
   REGISTERS_reg_7_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_7_2_port, QN => n_1307);
   REGISTERS_reg_7_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_7_1_port, QN => n_1308);
   REGISTERS_reg_7_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N295, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_7_0_port, QN => n_1309);
   REGISTERS_reg_8_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_8_31_port, QN => n_1310);
   REGISTERS_reg_8_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_8_30_port, QN => n_1311);
   REGISTERS_reg_8_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_8_29_port, QN => n_1312);
   REGISTERS_reg_8_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_8_28_port, QN => n_1313);
   REGISTERS_reg_8_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_8_27_port, QN => n_1314);
   REGISTERS_reg_8_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_8_26_port, QN => n_1315);
   REGISTERS_reg_8_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_8_25_port, QN => n_1316);
   REGISTERS_reg_8_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_8_24_port, QN => n_1317);
   REGISTERS_reg_8_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_8_23_port, QN => n_1318);
   REGISTERS_reg_8_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_8_22_port, QN => n_1319);
   REGISTERS_reg_8_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_8_21_port, QN => n_1320);
   REGISTERS_reg_8_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_8_20_port, QN => n_1321);
   REGISTERS_reg_8_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_8_19_port, QN => n_1322);
   REGISTERS_reg_8_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_8_18_port, QN => n_1323);
   REGISTERS_reg_8_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_8_17_port, QN => n_1324);
   REGISTERS_reg_8_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_8_16_port, QN => n_1325);
   REGISTERS_reg_8_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_8_15_port, QN => n_1326);
   REGISTERS_reg_8_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_8_14_port, QN => n_1327);
   REGISTERS_reg_8_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_8_13_port, QN => n_1328);
   REGISTERS_reg_8_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_8_12_port, QN => n_1329);
   REGISTERS_reg_8_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_8_11_port, QN => n_1330);
   REGISTERS_reg_8_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_8_10_port, QN => n_1331);
   REGISTERS_reg_8_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_8_9_port, QN => n_1332);
   REGISTERS_reg_8_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_8_8_port, QN => n_1333);
   REGISTERS_reg_8_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_8_7_port, QN => n_1334);
   REGISTERS_reg_8_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_8_6_port, QN => n_1335);
   REGISTERS_reg_8_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_8_5_port, QN => n_1336);
   REGISTERS_reg_8_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_8_4_port, QN => n_1337);
   REGISTERS_reg_8_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_8_3_port, QN => n_1338);
   REGISTERS_reg_8_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_8_2_port, QN => n_1339);
   REGISTERS_reg_8_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_8_1_port, QN => n_1340);
   REGISTERS_reg_8_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N294, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_8_0_port, QN => n_1341);
   REGISTERS_reg_9_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_9_31_port, QN => n_1342);
   REGISTERS_reg_9_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_9_30_port, QN => n_1343);
   REGISTERS_reg_9_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_9_29_port, QN => n_1344);
   REGISTERS_reg_9_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_9_28_port, QN => n_1345);
   REGISTERS_reg_9_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_9_27_port, QN => n_1346);
   REGISTERS_reg_9_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_9_26_port, QN => n_1347);
   REGISTERS_reg_9_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_9_25_port, QN => n_1348);
   REGISTERS_reg_9_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_9_24_port, QN => n_1349);
   REGISTERS_reg_9_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_9_23_port, QN => n_1350);
   REGISTERS_reg_9_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_9_22_port, QN => n_1351);
   REGISTERS_reg_9_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_9_21_port, QN => n_1352);
   REGISTERS_reg_9_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_9_20_port, QN => n_1353);
   REGISTERS_reg_9_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_9_19_port, QN => n_1354);
   REGISTERS_reg_9_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_9_18_port, QN => n_1355);
   REGISTERS_reg_9_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_9_17_port, QN => n_1356);
   REGISTERS_reg_9_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_9_16_port, QN => n_1357);
   REGISTERS_reg_9_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_9_15_port, QN => n_1358);
   REGISTERS_reg_9_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_9_14_port, QN => n_1359);
   REGISTERS_reg_9_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_9_13_port, QN => n_1360);
   REGISTERS_reg_9_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_9_12_port, QN => n_1361);
   REGISTERS_reg_9_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_9_11_port, QN => n_1362);
   REGISTERS_reg_9_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_9_10_port, QN => n_1363);
   REGISTERS_reg_9_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_9_9_port, QN => n_1364);
   REGISTERS_reg_9_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_9_8_port, QN => n_1365);
   REGISTERS_reg_9_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_9_7_port, QN => n_1366);
   REGISTERS_reg_9_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_9_6_port, QN => n_1367);
   REGISTERS_reg_9_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_9_5_port, QN => n_1368);
   REGISTERS_reg_9_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_9_4_port, QN => n_1369);
   REGISTERS_reg_9_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_9_3_port, QN => n_1370);
   REGISTERS_reg_9_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_9_2_port, QN => n_1371);
   REGISTERS_reg_9_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_9_1_port, QN => n_1372);
   REGISTERS_reg_9_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N293, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_9_0_port, QN => n_1373);
   REGISTERS_reg_10_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_10_31_port, QN => n_1374
               );
   REGISTERS_reg_10_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_10_30_port, QN => n_1375
               );
   REGISTERS_reg_10_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_10_29_port, QN => n_1376
               );
   REGISTERS_reg_10_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_10_28_port, QN => n_1377
               );
   REGISTERS_reg_10_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_10_27_port, QN => n_1378
               );
   REGISTERS_reg_10_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_10_26_port, QN => n_1379
               );
   REGISTERS_reg_10_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_10_25_port, QN => n_1380
               );
   REGISTERS_reg_10_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_10_24_port, QN => n_1381
               );
   REGISTERS_reg_10_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_10_23_port, QN => n_1382
               );
   REGISTERS_reg_10_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_10_22_port, QN => n_1383
               );
   REGISTERS_reg_10_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_10_21_port, QN => n_1384
               );
   REGISTERS_reg_10_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_10_20_port, QN => n_1385
               );
   REGISTERS_reg_10_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_10_19_port, QN => n_1386
               );
   REGISTERS_reg_10_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_10_18_port, QN => n_1387
               );
   REGISTERS_reg_10_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_10_17_port, QN => n_1388
               );
   REGISTERS_reg_10_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_10_16_port, QN => n_1389
               );
   REGISTERS_reg_10_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_10_15_port, QN => n_1390
               );
   REGISTERS_reg_10_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_10_14_port, QN => n_1391
               );
   REGISTERS_reg_10_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_10_13_port, QN => n_1392
               );
   REGISTERS_reg_10_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_10_12_port, QN => n_1393
               );
   REGISTERS_reg_10_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_10_11_port, QN => n_1394
               );
   REGISTERS_reg_10_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_10_10_port, QN => n_1395
               );
   REGISTERS_reg_10_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_10_9_port, QN => n_1396);
   REGISTERS_reg_10_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_10_8_port, QN => n_1397);
   REGISTERS_reg_10_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_10_7_port, QN => n_1398);
   REGISTERS_reg_10_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_10_6_port, QN => n_1399);
   REGISTERS_reg_10_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_10_5_port, QN => n_1400);
   REGISTERS_reg_10_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_10_4_port, QN => n_1401);
   REGISTERS_reg_10_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_10_3_port, QN => n_1402);
   REGISTERS_reg_10_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_10_2_port, QN => n_1403);
   REGISTERS_reg_10_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_10_1_port, QN => n_1404);
   REGISTERS_reg_10_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N292, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_10_0_port, QN => n_1405);
   REGISTERS_reg_11_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_11_31_port, QN => n_1406
               );
   REGISTERS_reg_11_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_11_30_port, QN => n_1407
               );
   REGISTERS_reg_11_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_11_29_port, QN => n_1408
               );
   REGISTERS_reg_11_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_11_28_port, QN => n_1409
               );
   REGISTERS_reg_11_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_11_27_port, QN => n_1410
               );
   REGISTERS_reg_11_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_11_26_port, QN => n_1411
               );
   REGISTERS_reg_11_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_11_25_port, QN => n_1412
               );
   REGISTERS_reg_11_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_11_24_port, QN => n_1413
               );
   REGISTERS_reg_11_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_11_23_port, QN => n_1414
               );
   REGISTERS_reg_11_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_11_22_port, QN => n_1415
               );
   REGISTERS_reg_11_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_11_21_port, QN => n_1416
               );
   REGISTERS_reg_11_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_11_20_port, QN => n_1417
               );
   REGISTERS_reg_11_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_11_19_port, QN => n_1418
               );
   REGISTERS_reg_11_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_11_18_port, QN => n_1419
               );
   REGISTERS_reg_11_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_11_17_port, QN => n_1420
               );
   REGISTERS_reg_11_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_11_16_port, QN => n_1421
               );
   REGISTERS_reg_11_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_11_15_port, QN => n_1422
               );
   REGISTERS_reg_11_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_11_14_port, QN => n_1423
               );
   REGISTERS_reg_11_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_11_13_port, QN => n_1424
               );
   REGISTERS_reg_11_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_11_12_port, QN => n_1425
               );
   REGISTERS_reg_11_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_11_11_port, QN => n_1426
               );
   REGISTERS_reg_11_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_11_10_port, QN => n_1427
               );
   REGISTERS_reg_11_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_11_9_port, QN => n_1428);
   REGISTERS_reg_11_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_11_8_port, QN => n_1429);
   REGISTERS_reg_11_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_11_7_port, QN => n_1430);
   REGISTERS_reg_11_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_11_6_port, QN => n_1431);
   REGISTERS_reg_11_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_11_5_port, QN => n_1432);
   REGISTERS_reg_11_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_11_4_port, QN => n_1433);
   REGISTERS_reg_11_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_11_3_port, QN => n_1434);
   REGISTERS_reg_11_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_11_2_port, QN => n_1435);
   REGISTERS_reg_11_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_11_1_port, QN => n_1436);
   REGISTERS_reg_11_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N291, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_11_0_port, QN => n_1437);
   REGISTERS_reg_12_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_12_31_port, QN => n_1438
               );
   REGISTERS_reg_12_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_12_30_port, QN => n_1439
               );
   REGISTERS_reg_12_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_12_29_port, QN => n_1440
               );
   REGISTERS_reg_12_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_12_28_port, QN => n_1441
               );
   REGISTERS_reg_12_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_12_27_port, QN => n_1442
               );
   REGISTERS_reg_12_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_12_26_port, QN => n_1443
               );
   REGISTERS_reg_12_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_12_25_port, QN => n_1444
               );
   REGISTERS_reg_12_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_12_24_port, QN => n_1445
               );
   REGISTERS_reg_12_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_12_23_port, QN => n_1446
               );
   REGISTERS_reg_12_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_12_22_port, QN => n_1447
               );
   REGISTERS_reg_12_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_12_21_port, QN => n_1448
               );
   REGISTERS_reg_12_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_12_20_port, QN => n_1449
               );
   REGISTERS_reg_12_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_12_19_port, QN => n_1450
               );
   REGISTERS_reg_12_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_12_18_port, QN => n_1451
               );
   REGISTERS_reg_12_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_12_17_port, QN => n_1452
               );
   REGISTERS_reg_12_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_12_16_port, QN => n_1453
               );
   REGISTERS_reg_12_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_12_15_port, QN => n_1454
               );
   REGISTERS_reg_12_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_12_14_port, QN => n_1455
               );
   REGISTERS_reg_12_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_12_13_port, QN => n_1456
               );
   REGISTERS_reg_12_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_12_12_port, QN => n_1457
               );
   REGISTERS_reg_12_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_12_11_port, QN => n_1458
               );
   REGISTERS_reg_12_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_12_10_port, QN => n_1459
               );
   REGISTERS_reg_12_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_12_9_port, QN => n_1460);
   REGISTERS_reg_12_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_12_8_port, QN => n_1461);
   REGISTERS_reg_12_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_12_7_port, QN => n_1462);
   REGISTERS_reg_12_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_12_6_port, QN => n_1463);
   REGISTERS_reg_12_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_12_5_port, QN => n_1464);
   REGISTERS_reg_12_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_12_4_port, QN => n_1465);
   REGISTERS_reg_12_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_12_3_port, QN => n_1466);
   REGISTERS_reg_12_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_12_2_port, QN => n_1467);
   REGISTERS_reg_12_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_12_1_port, QN => n_1468);
   REGISTERS_reg_12_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N290, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_12_0_port, QN => n_1469);
   REGISTERS_reg_13_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_13_31_port, QN => n_1470
               );
   REGISTERS_reg_13_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_13_30_port, QN => n_1471
               );
   REGISTERS_reg_13_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_13_29_port, QN => n_1472
               );
   REGISTERS_reg_13_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_13_28_port, QN => n_1473
               );
   REGISTERS_reg_13_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_13_27_port, QN => n_1474
               );
   REGISTERS_reg_13_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_13_26_port, QN => n_1475
               );
   REGISTERS_reg_13_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_13_25_port, QN => n_1476
               );
   REGISTERS_reg_13_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_13_24_port, QN => n_1477
               );
   REGISTERS_reg_13_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_13_23_port, QN => n_1478
               );
   REGISTERS_reg_13_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_13_22_port, QN => n_1479
               );
   REGISTERS_reg_13_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_13_21_port, QN => n_1480
               );
   REGISTERS_reg_13_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_13_20_port, QN => n_1481
               );
   REGISTERS_reg_13_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_13_19_port, QN => n_1482
               );
   REGISTERS_reg_13_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_13_18_port, QN => n_1483
               );
   REGISTERS_reg_13_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_13_17_port, QN => n_1484
               );
   REGISTERS_reg_13_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_13_16_port, QN => n_1485
               );
   REGISTERS_reg_13_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_13_15_port, QN => n_1486
               );
   REGISTERS_reg_13_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_13_14_port, QN => n_1487
               );
   REGISTERS_reg_13_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_13_13_port, QN => n_1488
               );
   REGISTERS_reg_13_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_13_12_port, QN => n_1489
               );
   REGISTERS_reg_13_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_13_11_port, QN => n_1490
               );
   REGISTERS_reg_13_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_13_10_port, QN => n_1491
               );
   REGISTERS_reg_13_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_13_9_port, QN => n_1492);
   REGISTERS_reg_13_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_13_8_port, QN => n_1493);
   REGISTERS_reg_13_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_13_7_port, QN => n_1494);
   REGISTERS_reg_13_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_13_6_port, QN => n_1495);
   REGISTERS_reg_13_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_13_5_port, QN => n_1496);
   REGISTERS_reg_13_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_13_4_port, QN => n_1497);
   REGISTERS_reg_13_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_13_3_port, QN => n_1498);
   REGISTERS_reg_13_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_13_2_port, QN => n_1499);
   REGISTERS_reg_13_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_13_1_port, QN => n_1500);
   REGISTERS_reg_13_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N289, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_13_0_port, QN => n_1501);
   REGISTERS_reg_14_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_14_31_port, QN => n_1502
               );
   REGISTERS_reg_14_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_14_30_port, QN => n_1503
               );
   REGISTERS_reg_14_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_14_29_port, QN => n_1504
               );
   REGISTERS_reg_14_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_14_28_port, QN => n_1505
               );
   REGISTERS_reg_14_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_14_27_port, QN => n_1506
               );
   REGISTERS_reg_14_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_14_26_port, QN => n_1507
               );
   REGISTERS_reg_14_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_14_25_port, QN => n_1508
               );
   REGISTERS_reg_14_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_14_24_port, QN => n_1509
               );
   REGISTERS_reg_14_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_14_23_port, QN => n_1510
               );
   REGISTERS_reg_14_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_14_22_port, QN => n_1511
               );
   REGISTERS_reg_14_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_14_21_port, QN => n_1512
               );
   REGISTERS_reg_14_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_14_20_port, QN => n_1513
               );
   REGISTERS_reg_14_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_14_19_port, QN => n_1514
               );
   REGISTERS_reg_14_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_14_18_port, QN => n_1515
               );
   REGISTERS_reg_14_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_14_17_port, QN => n_1516
               );
   REGISTERS_reg_14_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_14_16_port, QN => n_1517
               );
   REGISTERS_reg_14_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_14_15_port, QN => n_1518
               );
   REGISTERS_reg_14_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_14_14_port, QN => n_1519
               );
   REGISTERS_reg_14_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_14_13_port, QN => n_1520
               );
   REGISTERS_reg_14_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_14_12_port, QN => n_1521
               );
   REGISTERS_reg_14_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_14_11_port, QN => n_1522
               );
   REGISTERS_reg_14_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_14_10_port, QN => n_1523
               );
   REGISTERS_reg_14_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_14_9_port, QN => n_1524);
   REGISTERS_reg_14_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_14_8_port, QN => n_1525);
   REGISTERS_reg_14_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_14_7_port, QN => n_1526);
   REGISTERS_reg_14_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_14_6_port, QN => n_1527);
   REGISTERS_reg_14_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_14_5_port, QN => n_1528);
   REGISTERS_reg_14_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_14_4_port, QN => n_1529);
   REGISTERS_reg_14_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_14_3_port, QN => n_1530);
   REGISTERS_reg_14_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_14_2_port, QN => n_1531);
   REGISTERS_reg_14_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_14_1_port, QN => n_1532);
   REGISTERS_reg_14_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N288, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_14_0_port, QN => n_1533);
   REGISTERS_reg_15_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_15_31_port, QN => n_1534
               );
   REGISTERS_reg_15_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_15_30_port, QN => n_1535
               );
   REGISTERS_reg_15_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_15_29_port, QN => n_1536
               );
   REGISTERS_reg_15_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_15_28_port, QN => n_1537
               );
   REGISTERS_reg_15_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_15_27_port, QN => n_1538
               );
   REGISTERS_reg_15_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_15_26_port, QN => n_1539
               );
   REGISTERS_reg_15_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_15_25_port, QN => n_1540
               );
   REGISTERS_reg_15_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_15_24_port, QN => n_1541
               );
   REGISTERS_reg_15_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_15_23_port, QN => n_1542
               );
   REGISTERS_reg_15_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_15_22_port, QN => n_1543
               );
   REGISTERS_reg_15_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_15_21_port, QN => n_1544
               );
   REGISTERS_reg_15_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_15_20_port, QN => n_1545
               );
   REGISTERS_reg_15_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_15_19_port, QN => n_1546
               );
   REGISTERS_reg_15_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_15_18_port, QN => n_1547
               );
   REGISTERS_reg_15_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_15_17_port, QN => n_1548
               );
   REGISTERS_reg_15_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_15_16_port, QN => n_1549
               );
   REGISTERS_reg_15_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_15_15_port, QN => n_1550
               );
   REGISTERS_reg_15_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_15_14_port, QN => n_1551
               );
   REGISTERS_reg_15_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_15_13_port, QN => n_1552
               );
   REGISTERS_reg_15_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_15_12_port, QN => n_1553
               );
   REGISTERS_reg_15_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_15_11_port, QN => n_1554
               );
   REGISTERS_reg_15_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_15_10_port, QN => n_1555
               );
   REGISTERS_reg_15_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_15_9_port, QN => n_1556);
   REGISTERS_reg_15_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_15_8_port, QN => n_1557);
   REGISTERS_reg_15_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_15_7_port, QN => n_1558);
   REGISTERS_reg_15_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_15_6_port, QN => n_1559);
   REGISTERS_reg_15_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_15_5_port, QN => n_1560);
   REGISTERS_reg_15_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_15_4_port, QN => n_1561);
   REGISTERS_reg_15_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_15_3_port, QN => n_1562);
   REGISTERS_reg_15_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_15_2_port, QN => n_1563);
   REGISTERS_reg_15_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_15_1_port, QN => n_1564);
   REGISTERS_reg_15_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N287, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_15_0_port, QN => n_1565);
   REGISTERS_reg_16_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_16_31_port, QN => n_1566
               );
   REGISTERS_reg_16_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_16_30_port, QN => n_1567
               );
   REGISTERS_reg_16_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_16_29_port, QN => n_1568
               );
   REGISTERS_reg_16_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_16_28_port, QN => n_1569
               );
   REGISTERS_reg_16_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_16_27_port, QN => n_1570
               );
   REGISTERS_reg_16_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_16_26_port, QN => n_1571
               );
   REGISTERS_reg_16_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_16_25_port, QN => n_1572
               );
   REGISTERS_reg_16_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_16_24_port, QN => n_1573
               );
   REGISTERS_reg_16_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_16_23_port, QN => n_1574
               );
   REGISTERS_reg_16_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_16_22_port, QN => n_1575
               );
   REGISTERS_reg_16_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_16_21_port, QN => n_1576
               );
   REGISTERS_reg_16_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_16_20_port, QN => n_1577
               );
   REGISTERS_reg_16_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_16_19_port, QN => n_1578
               );
   REGISTERS_reg_16_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_16_18_port, QN => n_1579
               );
   REGISTERS_reg_16_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_16_17_port, QN => n_1580
               );
   REGISTERS_reg_16_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_16_16_port, QN => n_1581
               );
   REGISTERS_reg_16_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_16_15_port, QN => n_1582
               );
   REGISTERS_reg_16_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_16_14_port, QN => n_1583
               );
   REGISTERS_reg_16_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_16_13_port, QN => n_1584
               );
   REGISTERS_reg_16_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_16_12_port, QN => n_1585
               );
   REGISTERS_reg_16_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_16_11_port, QN => n_1586
               );
   REGISTERS_reg_16_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_16_10_port, QN => n_1587
               );
   REGISTERS_reg_16_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_16_9_port, QN => n_1588);
   REGISTERS_reg_16_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_16_8_port, QN => n_1589);
   REGISTERS_reg_16_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_16_7_port, QN => n_1590);
   REGISTERS_reg_16_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_16_6_port, QN => n_1591);
   REGISTERS_reg_16_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_16_5_port, QN => n_1592);
   REGISTERS_reg_16_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_16_4_port, QN => n_1593);
   REGISTERS_reg_16_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_16_3_port, QN => n_1594);
   REGISTERS_reg_16_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_16_2_port, QN => n_1595);
   REGISTERS_reg_16_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_16_1_port, QN => n_1596);
   REGISTERS_reg_16_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N286, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_16_0_port, QN => n_1597);
   REGISTERS_reg_17_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_17_31_port, QN => n_1598
               );
   REGISTERS_reg_17_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_17_30_port, QN => n_1599
               );
   REGISTERS_reg_17_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_17_29_port, QN => n_1600
               );
   REGISTERS_reg_17_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_17_28_port, QN => n_1601
               );
   REGISTERS_reg_17_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_17_27_port, QN => n_1602
               );
   REGISTERS_reg_17_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_17_26_port, QN => n_1603
               );
   REGISTERS_reg_17_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_17_25_port, QN => n_1604
               );
   REGISTERS_reg_17_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_17_24_port, QN => n_1605
               );
   REGISTERS_reg_17_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_17_23_port, QN => n_1606
               );
   REGISTERS_reg_17_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_17_22_port, QN => n_1607
               );
   REGISTERS_reg_17_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_17_21_port, QN => n_1608
               );
   REGISTERS_reg_17_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_17_20_port, QN => n_1609
               );
   REGISTERS_reg_17_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_17_19_port, QN => n_1610
               );
   REGISTERS_reg_17_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_17_18_port, QN => n_1611
               );
   REGISTERS_reg_17_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_17_17_port, QN => n_1612
               );
   REGISTERS_reg_17_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_17_16_port, QN => n_1613
               );
   REGISTERS_reg_17_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_17_15_port, QN => n_1614
               );
   REGISTERS_reg_17_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_17_14_port, QN => n_1615
               );
   REGISTERS_reg_17_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_17_13_port, QN => n_1616
               );
   REGISTERS_reg_17_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_17_12_port, QN => n_1617
               );
   REGISTERS_reg_17_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_17_11_port, QN => n_1618
               );
   REGISTERS_reg_17_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_17_10_port, QN => n_1619
               );
   REGISTERS_reg_17_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_17_9_port, QN => n_1620);
   REGISTERS_reg_17_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_17_8_port, QN => n_1621);
   REGISTERS_reg_17_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_17_7_port, QN => n_1622);
   REGISTERS_reg_17_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_17_6_port, QN => n_1623);
   REGISTERS_reg_17_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_17_5_port, QN => n_1624);
   REGISTERS_reg_17_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_17_4_port, QN => n_1625);
   REGISTERS_reg_17_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_17_3_port, QN => n_1626);
   REGISTERS_reg_17_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_17_2_port, QN => n_1627);
   REGISTERS_reg_17_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_17_1_port, QN => n_1628);
   REGISTERS_reg_17_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N285, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_17_0_port, QN => n_1629);
   REGISTERS_reg_18_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_18_31_port, QN => n_1630
               );
   REGISTERS_reg_18_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_18_30_port, QN => n_1631
               );
   REGISTERS_reg_18_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_18_29_port, QN => n_1632
               );
   REGISTERS_reg_18_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_18_28_port, QN => n_1633
               );
   REGISTERS_reg_18_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_18_27_port, QN => n_1634
               );
   REGISTERS_reg_18_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_18_26_port, QN => n_1635
               );
   REGISTERS_reg_18_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_18_25_port, QN => n_1636
               );
   REGISTERS_reg_18_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_18_24_port, QN => n_1637
               );
   REGISTERS_reg_18_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_18_23_port, QN => n_1638
               );
   REGISTERS_reg_18_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_18_22_port, QN => n_1639
               );
   REGISTERS_reg_18_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_18_21_port, QN => n_1640
               );
   REGISTERS_reg_18_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_18_20_port, QN => n_1641
               );
   REGISTERS_reg_18_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_18_19_port, QN => n_1642
               );
   REGISTERS_reg_18_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_18_18_port, QN => n_1643
               );
   REGISTERS_reg_18_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_18_17_port, QN => n_1644
               );
   REGISTERS_reg_18_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_18_16_port, QN => n_1645
               );
   REGISTERS_reg_18_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_18_15_port, QN => n_1646
               );
   REGISTERS_reg_18_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_18_14_port, QN => n_1647
               );
   REGISTERS_reg_18_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_18_13_port, QN => n_1648
               );
   REGISTERS_reg_18_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_18_12_port, QN => n_1649
               );
   REGISTERS_reg_18_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_18_11_port, QN => n_1650
               );
   REGISTERS_reg_18_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_18_10_port, QN => n_1651
               );
   REGISTERS_reg_18_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_18_9_port, QN => n_1652);
   REGISTERS_reg_18_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_18_8_port, QN => n_1653);
   REGISTERS_reg_18_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_18_7_port, QN => n_1654);
   REGISTERS_reg_18_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_18_6_port, QN => n_1655);
   REGISTERS_reg_18_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_18_5_port, QN => n_1656);
   REGISTERS_reg_18_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_18_4_port, QN => n_1657);
   REGISTERS_reg_18_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_18_3_port, QN => n_1658);
   REGISTERS_reg_18_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_18_2_port, QN => n_1659);
   REGISTERS_reg_18_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_18_1_port, QN => n_1660);
   REGISTERS_reg_18_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N284, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_18_0_port, QN => n_1661);
   REGISTERS_reg_19_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_19_31_port, QN => n_1662
               );
   REGISTERS_reg_19_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_19_30_port, QN => n_1663
               );
   REGISTERS_reg_19_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_19_29_port, QN => n_1664
               );
   REGISTERS_reg_19_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_19_28_port, QN => n_1665
               );
   REGISTERS_reg_19_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_19_27_port, QN => n_1666
               );
   REGISTERS_reg_19_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_19_26_port, QN => n_1667
               );
   REGISTERS_reg_19_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_19_25_port, QN => n_1668
               );
   REGISTERS_reg_19_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_19_24_port, QN => n_1669
               );
   REGISTERS_reg_19_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_19_23_port, QN => n_1670
               );
   REGISTERS_reg_19_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_19_22_port, QN => n_1671
               );
   REGISTERS_reg_19_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_19_21_port, QN => n_1672
               );
   REGISTERS_reg_19_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_19_20_port, QN => n_1673
               );
   REGISTERS_reg_19_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_19_19_port, QN => n_1674
               );
   REGISTERS_reg_19_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_19_18_port, QN => n_1675
               );
   REGISTERS_reg_19_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_19_17_port, QN => n_1676
               );
   REGISTERS_reg_19_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_19_16_port, QN => n_1677
               );
   REGISTERS_reg_19_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_19_15_port, QN => n_1678
               );
   REGISTERS_reg_19_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_19_14_port, QN => n_1679
               );
   REGISTERS_reg_19_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_19_13_port, QN => n_1680
               );
   REGISTERS_reg_19_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_19_12_port, QN => n_1681
               );
   REGISTERS_reg_19_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_19_11_port, QN => n_1682
               );
   REGISTERS_reg_19_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_19_10_port, QN => n_1683
               );
   REGISTERS_reg_19_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_19_9_port, QN => n_1684);
   REGISTERS_reg_19_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_19_8_port, QN => n_1685);
   REGISTERS_reg_19_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_19_7_port, QN => n_1686);
   REGISTERS_reg_19_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_19_6_port, QN => n_1687);
   REGISTERS_reg_19_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_19_5_port, QN => n_1688);
   REGISTERS_reg_19_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_19_4_port, QN => n_1689);
   REGISTERS_reg_19_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_19_3_port, QN => n_1690);
   REGISTERS_reg_19_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_19_2_port, QN => n_1691);
   REGISTERS_reg_19_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_19_1_port, QN => n_1692);
   REGISTERS_reg_19_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N283, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_19_0_port, QN => n_1693);
   REGISTERS_reg_20_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_20_31_port, QN => n_1694
               );
   REGISTERS_reg_20_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_20_30_port, QN => n_1695
               );
   REGISTERS_reg_20_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_20_29_port, QN => n_1696
               );
   REGISTERS_reg_20_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_20_28_port, QN => n_1697
               );
   REGISTERS_reg_20_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_20_27_port, QN => n_1698
               );
   REGISTERS_reg_20_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_20_26_port, QN => n_1699
               );
   REGISTERS_reg_20_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_20_25_port, QN => n_1700
               );
   REGISTERS_reg_20_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_20_24_port, QN => n_1701
               );
   REGISTERS_reg_20_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_20_23_port, QN => n_1702
               );
   REGISTERS_reg_20_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_20_22_port, QN => n_1703
               );
   REGISTERS_reg_20_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_20_21_port, QN => n_1704
               );
   REGISTERS_reg_20_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_20_20_port, QN => n_1705
               );
   REGISTERS_reg_20_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_20_19_port, QN => n_1706
               );
   REGISTERS_reg_20_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_20_18_port, QN => n_1707
               );
   REGISTERS_reg_20_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_20_17_port, QN => n_1708
               );
   REGISTERS_reg_20_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_20_16_port, QN => n_1709
               );
   REGISTERS_reg_20_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_20_15_port, QN => n_1710
               );
   REGISTERS_reg_20_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_20_14_port, QN => n_1711
               );
   REGISTERS_reg_20_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_20_13_port, QN => n_1712
               );
   REGISTERS_reg_20_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_20_12_port, QN => n_1713
               );
   REGISTERS_reg_20_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_20_11_port, QN => n_1714
               );
   REGISTERS_reg_20_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_20_10_port, QN => n_1715
               );
   REGISTERS_reg_20_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_20_9_port, QN => n_1716);
   REGISTERS_reg_20_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_20_8_port, QN => n_1717);
   REGISTERS_reg_20_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_20_7_port, QN => n_1718);
   REGISTERS_reg_20_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_20_6_port, QN => n_1719);
   REGISTERS_reg_20_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_20_5_port, QN => n_1720);
   REGISTERS_reg_20_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_20_4_port, QN => n_1721);
   REGISTERS_reg_20_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_20_3_port, QN => n_1722);
   REGISTERS_reg_20_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_20_2_port, QN => n_1723);
   REGISTERS_reg_20_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_20_1_port, QN => n_1724);
   REGISTERS_reg_20_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N282, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_20_0_port, QN => n_1725);
   REGISTERS_reg_21_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_21_31_port, QN => n_1726
               );
   REGISTERS_reg_21_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_21_30_port, QN => n_1727
               );
   REGISTERS_reg_21_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_21_29_port, QN => n_1728
               );
   REGISTERS_reg_21_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_21_28_port, QN => n_1729
               );
   REGISTERS_reg_21_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_21_27_port, QN => n_1730
               );
   REGISTERS_reg_21_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_21_26_port, QN => n_1731
               );
   REGISTERS_reg_21_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_21_25_port, QN => n_1732
               );
   REGISTERS_reg_21_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_21_24_port, QN => n_1733
               );
   REGISTERS_reg_21_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_21_23_port, QN => n_1734
               );
   REGISTERS_reg_21_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_21_22_port, QN => n_1735
               );
   REGISTERS_reg_21_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_21_21_port, QN => n_1736
               );
   REGISTERS_reg_21_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_21_20_port, QN => n_1737
               );
   REGISTERS_reg_21_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_21_19_port, QN => n_1738
               );
   REGISTERS_reg_21_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_21_18_port, QN => n_1739
               );
   REGISTERS_reg_21_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_21_17_port, QN => n_1740
               );
   REGISTERS_reg_21_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_21_16_port, QN => n_1741
               );
   REGISTERS_reg_21_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_21_15_port, QN => n_1742
               );
   REGISTERS_reg_21_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_21_14_port, QN => n_1743
               );
   REGISTERS_reg_21_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_21_13_port, QN => n_1744
               );
   REGISTERS_reg_21_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_21_12_port, QN => n_1745
               );
   REGISTERS_reg_21_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_21_11_port, QN => n_1746
               );
   REGISTERS_reg_21_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_21_10_port, QN => n_1747
               );
   REGISTERS_reg_21_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_21_9_port, QN => n_1748);
   REGISTERS_reg_21_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_21_8_port, QN => n_1749);
   REGISTERS_reg_21_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_21_7_port, QN => n_1750);
   REGISTERS_reg_21_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_21_6_port, QN => n_1751);
   REGISTERS_reg_21_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_21_5_port, QN => n_1752);
   REGISTERS_reg_21_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_21_4_port, QN => n_1753);
   REGISTERS_reg_21_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_21_3_port, QN => n_1754);
   REGISTERS_reg_21_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_21_2_port, QN => n_1755);
   REGISTERS_reg_21_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_21_1_port, QN => n_1756);
   REGISTERS_reg_21_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N281, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_21_0_port, QN => n_1757);
   REGISTERS_reg_22_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_22_31_port, QN => n_1758
               );
   REGISTERS_reg_22_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_22_30_port, QN => n_1759
               );
   REGISTERS_reg_22_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_22_29_port, QN => n_1760
               );
   REGISTERS_reg_22_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_22_28_port, QN => n_1761
               );
   REGISTERS_reg_22_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_22_27_port, QN => n_1762
               );
   REGISTERS_reg_22_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_22_26_port, QN => n_1763
               );
   REGISTERS_reg_22_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_22_25_port, QN => n_1764
               );
   REGISTERS_reg_22_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_22_24_port, QN => n_1765
               );
   REGISTERS_reg_22_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_22_23_port, QN => n_1766
               );
   REGISTERS_reg_22_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_22_22_port, QN => n_1767
               );
   REGISTERS_reg_22_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_22_21_port, QN => n_1768
               );
   REGISTERS_reg_22_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_22_20_port, QN => n_1769
               );
   REGISTERS_reg_22_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_22_19_port, QN => n_1770
               );
   REGISTERS_reg_22_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_22_18_port, QN => n_1771
               );
   REGISTERS_reg_22_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_22_17_port, QN => n_1772
               );
   REGISTERS_reg_22_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_22_16_port, QN => n_1773
               );
   REGISTERS_reg_22_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_22_15_port, QN => n_1774
               );
   REGISTERS_reg_22_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_22_14_port, QN => n_1775
               );
   REGISTERS_reg_22_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_22_13_port, QN => n_1776
               );
   REGISTERS_reg_22_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_22_12_port, QN => n_1777
               );
   REGISTERS_reg_22_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_22_11_port, QN => n_1778
               );
   REGISTERS_reg_22_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_22_10_port, QN => n_1779
               );
   REGISTERS_reg_22_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_22_9_port, QN => n_1780);
   REGISTERS_reg_22_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_22_8_port, QN => n_1781);
   REGISTERS_reg_22_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_22_7_port, QN => n_1782);
   REGISTERS_reg_22_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_22_6_port, QN => n_1783);
   REGISTERS_reg_22_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_22_5_port, QN => n_1784);
   REGISTERS_reg_22_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_22_4_port, QN => n_1785);
   REGISTERS_reg_22_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_22_3_port, QN => n_1786);
   REGISTERS_reg_22_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_22_2_port, QN => n_1787);
   REGISTERS_reg_22_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_22_1_port, QN => n_1788);
   REGISTERS_reg_22_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N280, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_22_0_port, QN => n_1789);
   REGISTERS_reg_23_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_23_31_port, QN => n_1790
               );
   REGISTERS_reg_23_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_23_30_port, QN => n_1791
               );
   REGISTERS_reg_23_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_23_29_port, QN => n_1792
               );
   REGISTERS_reg_23_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_23_28_port, QN => n_1793
               );
   REGISTERS_reg_23_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_23_27_port, QN => n_1794
               );
   REGISTERS_reg_23_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_23_26_port, QN => n_1795
               );
   REGISTERS_reg_23_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_23_25_port, QN => n_1796
               );
   REGISTERS_reg_23_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_23_24_port, QN => n_1797
               );
   REGISTERS_reg_23_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_23_23_port, QN => n_1798
               );
   REGISTERS_reg_23_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_23_22_port, QN => n_1799
               );
   REGISTERS_reg_23_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_23_21_port, QN => n_1800
               );
   REGISTERS_reg_23_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_23_20_port, QN => n_1801
               );
   REGISTERS_reg_23_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_23_19_port, QN => n_1802
               );
   REGISTERS_reg_23_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_23_18_port, QN => n_1803
               );
   REGISTERS_reg_23_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_23_17_port, QN => n_1804
               );
   REGISTERS_reg_23_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_23_16_port, QN => n_1805
               );
   REGISTERS_reg_23_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_23_15_port, QN => n_1806
               );
   REGISTERS_reg_23_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_23_14_port, QN => n_1807
               );
   REGISTERS_reg_23_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_23_13_port, QN => n_1808
               );
   REGISTERS_reg_23_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_23_12_port, QN => n_1809
               );
   REGISTERS_reg_23_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_23_11_port, QN => n_1810
               );
   REGISTERS_reg_23_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_23_10_port, QN => n_1811
               );
   REGISTERS_reg_23_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_23_9_port, QN => n_1812);
   REGISTERS_reg_23_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_23_8_port, QN => n_1813);
   REGISTERS_reg_23_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_23_7_port, QN => n_1814);
   REGISTERS_reg_23_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_23_6_port, QN => n_1815);
   REGISTERS_reg_23_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_23_5_port, QN => n_1816);
   REGISTERS_reg_23_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_23_4_port, QN => n_1817);
   REGISTERS_reg_23_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_23_3_port, QN => n_1818);
   REGISTERS_reg_23_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_23_2_port, QN => n_1819);
   REGISTERS_reg_23_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_23_1_port, QN => n_1820);
   REGISTERS_reg_23_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N279, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_23_0_port, QN => n_1821);
   REGISTERS_reg_24_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_24_31_port, QN => n_1822
               );
   REGISTERS_reg_24_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_24_30_port, QN => n_1823
               );
   REGISTERS_reg_24_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_24_29_port, QN => n_1824
               );
   REGISTERS_reg_24_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_24_28_port, QN => n_1825
               );
   REGISTERS_reg_24_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_24_27_port, QN => n_1826
               );
   REGISTERS_reg_24_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_24_26_port, QN => n_1827
               );
   REGISTERS_reg_24_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_24_25_port, QN => n_1828
               );
   REGISTERS_reg_24_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_24_24_port, QN => n_1829
               );
   REGISTERS_reg_24_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_24_23_port, QN => n_1830
               );
   REGISTERS_reg_24_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_24_22_port, QN => n_1831
               );
   REGISTERS_reg_24_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_24_21_port, QN => n_1832
               );
   REGISTERS_reg_24_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_24_20_port, QN => n_1833
               );
   REGISTERS_reg_24_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_24_19_port, QN => n_1834
               );
   REGISTERS_reg_24_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_24_18_port, QN => n_1835
               );
   REGISTERS_reg_24_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_24_17_port, QN => n_1836
               );
   REGISTERS_reg_24_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_24_16_port, QN => n_1837
               );
   REGISTERS_reg_24_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_24_15_port, QN => n_1838
               );
   REGISTERS_reg_24_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_24_14_port, QN => n_1839
               );
   REGISTERS_reg_24_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_24_13_port, QN => n_1840
               );
   REGISTERS_reg_24_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_24_12_port, QN => n_1841
               );
   REGISTERS_reg_24_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_24_11_port, QN => n_1842
               );
   REGISTERS_reg_24_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_24_10_port, QN => n_1843
               );
   REGISTERS_reg_24_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_24_9_port, QN => n_1844);
   REGISTERS_reg_24_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_24_8_port, QN => n_1845);
   REGISTERS_reg_24_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_24_7_port, QN => n_1846);
   REGISTERS_reg_24_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_24_6_port, QN => n_1847);
   REGISTERS_reg_24_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_24_5_port, QN => n_1848);
   REGISTERS_reg_24_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_24_4_port, QN => n_1849);
   REGISTERS_reg_24_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_24_3_port, QN => n_1850);
   REGISTERS_reg_24_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_24_2_port, QN => n_1851);
   REGISTERS_reg_24_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_24_1_port, QN => n_1852);
   REGISTERS_reg_24_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N278, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_24_0_port, QN => n_1853);
   REGISTERS_reg_25_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_25_31_port, QN => n_1854
               );
   REGISTERS_reg_25_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_25_30_port, QN => n_1855
               );
   REGISTERS_reg_25_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_25_29_port, QN => n_1856
               );
   REGISTERS_reg_25_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_25_28_port, QN => n_1857
               );
   REGISTERS_reg_25_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_25_27_port, QN => n_1858
               );
   REGISTERS_reg_25_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_25_26_port, QN => n_1859
               );
   REGISTERS_reg_25_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_25_25_port, QN => n_1860
               );
   REGISTERS_reg_25_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_25_24_port, QN => n_1861
               );
   REGISTERS_reg_25_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_25_23_port, QN => n_1862
               );
   REGISTERS_reg_25_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_25_22_port, QN => n_1863
               );
   REGISTERS_reg_25_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_25_21_port, QN => n_1864
               );
   REGISTERS_reg_25_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_25_20_port, QN => n_1865
               );
   REGISTERS_reg_25_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_25_19_port, QN => n_1866
               );
   REGISTERS_reg_25_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_25_18_port, QN => n_1867
               );
   REGISTERS_reg_25_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_25_17_port, QN => n_1868
               );
   REGISTERS_reg_25_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_25_16_port, QN => n_1869
               );
   REGISTERS_reg_25_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_25_15_port, QN => n_1870
               );
   REGISTERS_reg_25_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_25_14_port, QN => n_1871
               );
   REGISTERS_reg_25_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_25_13_port, QN => n_1872
               );
   REGISTERS_reg_25_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_25_12_port, QN => n_1873
               );
   REGISTERS_reg_25_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_25_11_port, QN => n_1874
               );
   REGISTERS_reg_25_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_25_10_port, QN => n_1875
               );
   REGISTERS_reg_25_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_25_9_port, QN => n_1876);
   REGISTERS_reg_25_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_25_8_port, QN => n_1877);
   REGISTERS_reg_25_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_25_7_port, QN => n_1878);
   REGISTERS_reg_25_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_25_6_port, QN => n_1879);
   REGISTERS_reg_25_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_25_5_port, QN => n_1880);
   REGISTERS_reg_25_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_25_4_port, QN => n_1881);
   REGISTERS_reg_25_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_25_3_port, QN => n_1882);
   REGISTERS_reg_25_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_25_2_port, QN => n_1883);
   REGISTERS_reg_25_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_25_1_port, QN => n_1884);
   REGISTERS_reg_25_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N277, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_25_0_port, QN => n_1885);
   REGISTERS_reg_26_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_26_31_port, QN => n_1886
               );
   REGISTERS_reg_26_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_26_30_port, QN => n_1887
               );
   REGISTERS_reg_26_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_26_29_port, QN => n_1888
               );
   REGISTERS_reg_26_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_26_28_port, QN => n_1889
               );
   REGISTERS_reg_26_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_26_27_port, QN => n_1890
               );
   REGISTERS_reg_26_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_26_26_port, QN => n_1891
               );
   REGISTERS_reg_26_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_26_25_port, QN => n_1892
               );
   REGISTERS_reg_26_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_26_24_port, QN => n_1893
               );
   REGISTERS_reg_26_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_26_23_port, QN => n_1894
               );
   REGISTERS_reg_26_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_26_22_port, QN => n_1895
               );
   REGISTERS_reg_26_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_26_21_port, QN => n_1896
               );
   REGISTERS_reg_26_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_26_20_port, QN => n_1897
               );
   REGISTERS_reg_26_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_26_19_port, QN => n_1898
               );
   REGISTERS_reg_26_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_26_18_port, QN => n_1899
               );
   REGISTERS_reg_26_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_26_17_port, QN => n_1900
               );
   REGISTERS_reg_26_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_26_16_port, QN => n_1901
               );
   REGISTERS_reg_26_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_26_15_port, QN => n_1902
               );
   REGISTERS_reg_26_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_26_14_port, QN => n_1903
               );
   REGISTERS_reg_26_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_26_13_port, QN => n_1904
               );
   REGISTERS_reg_26_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_26_12_port, QN => n_1905
               );
   REGISTERS_reg_26_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_26_11_port, QN => n_1906
               );
   REGISTERS_reg_26_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_26_10_port, QN => n_1907
               );
   REGISTERS_reg_26_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_26_9_port, QN => n_1908);
   REGISTERS_reg_26_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_26_8_port, QN => n_1909);
   REGISTERS_reg_26_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_26_7_port, QN => n_1910);
   REGISTERS_reg_26_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_26_6_port, QN => n_1911);
   REGISTERS_reg_26_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_26_5_port, QN => n_1912);
   REGISTERS_reg_26_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_26_4_port, QN => n_1913);
   REGISTERS_reg_26_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_26_3_port, QN => n_1914);
   REGISTERS_reg_26_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_26_2_port, QN => n_1915);
   REGISTERS_reg_26_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_26_1_port, QN => n_1916);
   REGISTERS_reg_26_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N276, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_26_0_port, QN => n_1917);
   REGISTERS_reg_27_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_27_31_port, QN => n_1918
               );
   REGISTERS_reg_27_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_27_30_port, QN => n_1919
               );
   REGISTERS_reg_27_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_27_29_port, QN => n_1920
               );
   REGISTERS_reg_27_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_27_28_port, QN => n_1921
               );
   REGISTERS_reg_27_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_27_27_port, QN => n_1922
               );
   REGISTERS_reg_27_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_27_26_port, QN => n_1923
               );
   REGISTERS_reg_27_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_27_25_port, QN => n_1924
               );
   REGISTERS_reg_27_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_27_24_port, QN => n_1925
               );
   REGISTERS_reg_27_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_27_23_port, QN => n_1926
               );
   REGISTERS_reg_27_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_27_22_port, QN => n_1927
               );
   REGISTERS_reg_27_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_27_21_port, QN => n_1928
               );
   REGISTERS_reg_27_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_27_20_port, QN => n_1929
               );
   REGISTERS_reg_27_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_27_19_port, QN => n_1930
               );
   REGISTERS_reg_27_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_27_18_port, QN => n_1931
               );
   REGISTERS_reg_27_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_27_17_port, QN => n_1932
               );
   REGISTERS_reg_27_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_27_16_port, QN => n_1933
               );
   REGISTERS_reg_27_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_27_15_port, QN => n_1934
               );
   REGISTERS_reg_27_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_27_14_port, QN => n_1935
               );
   REGISTERS_reg_27_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_27_13_port, QN => n_1936
               );
   REGISTERS_reg_27_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_27_12_port, QN => n_1937
               );
   REGISTERS_reg_27_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_27_11_port, QN => n_1938
               );
   REGISTERS_reg_27_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_27_10_port, QN => n_1939
               );
   REGISTERS_reg_27_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_27_9_port, QN => n_1940);
   REGISTERS_reg_27_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_27_8_port, QN => n_1941);
   REGISTERS_reg_27_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_27_7_port, QN => n_1942);
   REGISTERS_reg_27_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_27_6_port, QN => n_1943);
   REGISTERS_reg_27_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_27_5_port, QN => n_1944);
   REGISTERS_reg_27_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_27_4_port, QN => n_1945);
   REGISTERS_reg_27_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_27_3_port, QN => n_1946);
   REGISTERS_reg_27_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_27_2_port, QN => n_1947);
   REGISTERS_reg_27_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_27_1_port, QN => n_1948);
   REGISTERS_reg_27_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N275, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_27_0_port, QN => n_1949);
   REGISTERS_reg_28_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_28_31_port, QN => n_1950
               );
   REGISTERS_reg_28_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_28_30_port, QN => n_1951
               );
   REGISTERS_reg_28_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_28_29_port, QN => n_1952
               );
   REGISTERS_reg_28_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_28_28_port, QN => n_1953
               );
   REGISTERS_reg_28_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_28_27_port, QN => n_1954
               );
   REGISTERS_reg_28_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_28_26_port, QN => n_1955
               );
   REGISTERS_reg_28_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_28_25_port, QN => n_1956
               );
   REGISTERS_reg_28_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_28_24_port, QN => n_1957
               );
   REGISTERS_reg_28_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_28_23_port, QN => n_1958
               );
   REGISTERS_reg_28_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_28_22_port, QN => n_1959
               );
   REGISTERS_reg_28_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_28_21_port, QN => n_1960
               );
   REGISTERS_reg_28_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_28_20_port, QN => n_1961
               );
   REGISTERS_reg_28_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_28_19_port, QN => n_1962
               );
   REGISTERS_reg_28_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_28_18_port, QN => n_1963
               );
   REGISTERS_reg_28_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_28_17_port, QN => n_1964
               );
   REGISTERS_reg_28_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_28_16_port, QN => n_1965
               );
   REGISTERS_reg_28_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_28_15_port, QN => n_1966
               );
   REGISTERS_reg_28_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_28_14_port, QN => n_1967
               );
   REGISTERS_reg_28_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_28_13_port, QN => n_1968
               );
   REGISTERS_reg_28_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_28_12_port, QN => n_1969
               );
   REGISTERS_reg_28_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_28_11_port, QN => n_1970
               );
   REGISTERS_reg_28_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_28_10_port, QN => n_1971
               );
   REGISTERS_reg_28_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_28_9_port, QN => n_1972);
   REGISTERS_reg_28_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_28_8_port, QN => n_1973);
   REGISTERS_reg_28_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_28_7_port, QN => n_1974);
   REGISTERS_reg_28_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_28_6_port, QN => n_1975);
   REGISTERS_reg_28_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_28_5_port, QN => n_1976);
   REGISTERS_reg_28_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_28_4_port, QN => n_1977);
   REGISTERS_reg_28_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_28_3_port, QN => n_1978);
   REGISTERS_reg_28_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_28_2_port, QN => n_1979);
   REGISTERS_reg_28_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_28_1_port, QN => n_1980);
   REGISTERS_reg_28_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N274, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_28_0_port, QN => n_1981);
   REGISTERS_reg_29_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_29_31_port, QN => n_1982
               );
   REGISTERS_reg_29_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_29_30_port, QN => n_1983
               );
   REGISTERS_reg_29_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_29_29_port, QN => n_1984
               );
   REGISTERS_reg_29_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_29_28_port, QN => n_1985
               );
   REGISTERS_reg_29_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_29_27_port, QN => n_1986
               );
   REGISTERS_reg_29_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_29_26_port, QN => n_1987
               );
   REGISTERS_reg_29_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_29_25_port, QN => n_1988
               );
   REGISTERS_reg_29_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_29_24_port, QN => n_1989
               );
   REGISTERS_reg_29_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_29_23_port, QN => n_1990
               );
   REGISTERS_reg_29_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_29_22_port, QN => n_1991
               );
   REGISTERS_reg_29_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_29_21_port, QN => n_1992
               );
   REGISTERS_reg_29_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_29_20_port, QN => n_1993
               );
   REGISTERS_reg_29_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_29_19_port, QN => n_1994
               );
   REGISTERS_reg_29_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_29_18_port, QN => n_1995
               );
   REGISTERS_reg_29_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_29_17_port, QN => n_1996
               );
   REGISTERS_reg_29_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_29_16_port, QN => n_1997
               );
   REGISTERS_reg_29_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_29_15_port, QN => n_1998
               );
   REGISTERS_reg_29_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_29_14_port, QN => n_1999
               );
   REGISTERS_reg_29_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_29_13_port, QN => n_2000
               );
   REGISTERS_reg_29_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_29_12_port, QN => n_2001
               );
   REGISTERS_reg_29_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_29_11_port, QN => n_2002
               );
   REGISTERS_reg_29_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_29_10_port, QN => n_2003
               );
   REGISTERS_reg_29_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_29_9_port, QN => n_2004);
   REGISTERS_reg_29_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_29_8_port, QN => n_2005);
   REGISTERS_reg_29_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_29_7_port, QN => n_2006);
   REGISTERS_reg_29_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_29_6_port, QN => n_2007);
   REGISTERS_reg_29_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_29_5_port, QN => n_2008);
   REGISTERS_reg_29_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_29_4_port, QN => n_2009);
   REGISTERS_reg_29_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_29_3_port, QN => n_2010);
   REGISTERS_reg_29_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_29_2_port, QN => n_2011);
   REGISTERS_reg_29_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_29_1_port, QN => n_2012);
   REGISTERS_reg_29_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N273, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_29_0_port, QN => n_2013);
   REGISTERS_reg_30_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_30_31_port, QN => n_2014
               );
   REGISTERS_reg_30_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_30_30_port, QN => n_2015
               );
   REGISTERS_reg_30_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_30_29_port, QN => n_2016
               );
   REGISTERS_reg_30_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_30_28_port, QN => n_2017
               );
   REGISTERS_reg_30_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_30_27_port, QN => n_2018
               );
   REGISTERS_reg_30_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_30_26_port, QN => n_2019
               );
   REGISTERS_reg_30_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_30_25_port, QN => n_2020
               );
   REGISTERS_reg_30_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_30_24_port, QN => n_2021
               );
   REGISTERS_reg_30_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_30_23_port, QN => n_2022
               );
   REGISTERS_reg_30_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_30_22_port, QN => n_2023
               );
   REGISTERS_reg_30_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_30_21_port, QN => n_2024
               );
   REGISTERS_reg_30_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_30_20_port, QN => n_2025
               );
   REGISTERS_reg_30_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_30_19_port, QN => n_2026
               );
   REGISTERS_reg_30_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_30_18_port, QN => n_2027
               );
   REGISTERS_reg_30_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_30_17_port, QN => n_2028
               );
   REGISTERS_reg_30_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_30_16_port, QN => n_2029
               );
   REGISTERS_reg_30_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_30_15_port, QN => n_2030
               );
   REGISTERS_reg_30_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_30_14_port, QN => n_2031
               );
   REGISTERS_reg_30_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_30_13_port, QN => n_2032
               );
   REGISTERS_reg_30_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_30_12_port, QN => n_2033
               );
   REGISTERS_reg_30_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_30_11_port, QN => n_2034
               );
   REGISTERS_reg_30_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_30_10_port, QN => n_2035
               );
   REGISTERS_reg_30_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_30_9_port, QN => n_2036);
   REGISTERS_reg_30_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_30_8_port, QN => n_2037);
   REGISTERS_reg_30_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_30_7_port, QN => n_2038);
   REGISTERS_reg_30_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_30_6_port, QN => n_2039);
   REGISTERS_reg_30_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_30_5_port, QN => n_2040);
   REGISTERS_reg_30_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_30_4_port, QN => n_2041);
   REGISTERS_reg_30_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_30_3_port, QN => n_2042);
   REGISTERS_reg_30_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_30_2_port, QN => n_2043);
   REGISTERS_reg_30_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_30_1_port, QN => n_2044);
   REGISTERS_reg_30_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N272, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_30_0_port, QN => n_2045);
   REGISTERS_reg_31_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N271, 
               clocked_on => CLK_port, Q => REGISTERS_31_31_port, QN => n_2046
               );
   REGISTERS_reg_31_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N270, 
               clocked_on => CLK_port, Q => REGISTERS_31_30_port, QN => n_2047
               );
   REGISTERS_reg_31_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N269, 
               clocked_on => CLK_port, Q => REGISTERS_31_29_port, QN => n_2048
               );
   REGISTERS_reg_31_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N268, 
               clocked_on => CLK_port, Q => REGISTERS_31_28_port, QN => n_2049
               );
   REGISTERS_reg_31_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N267, 
               clocked_on => CLK_port, Q => REGISTERS_31_27_port, QN => n_2050
               );
   REGISTERS_reg_31_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N266, 
               clocked_on => CLK_port, Q => REGISTERS_31_26_port, QN => n_2051
               );
   REGISTERS_reg_31_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N265, 
               clocked_on => CLK_port, Q => REGISTERS_31_25_port, QN => n_2052
               );
   REGISTERS_reg_31_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N264, 
               clocked_on => CLK_port, Q => REGISTERS_31_24_port, QN => n_2053
               );
   REGISTERS_reg_31_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N263, 
               clocked_on => CLK_port, Q => REGISTERS_31_23_port, QN => n_2054
               );
   REGISTERS_reg_31_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N262, 
               clocked_on => CLK_port, Q => REGISTERS_31_22_port, QN => n_2055
               );
   REGISTERS_reg_31_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N261, 
               clocked_on => CLK_port, Q => REGISTERS_31_21_port, QN => n_2056
               );
   REGISTERS_reg_31_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N260, 
               clocked_on => CLK_port, Q => REGISTERS_31_20_port, QN => n_2057
               );
   REGISTERS_reg_31_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N259, 
               clocked_on => CLK_port, Q => REGISTERS_31_19_port, QN => n_2058
               );
   REGISTERS_reg_31_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N258, 
               clocked_on => CLK_port, Q => REGISTERS_31_18_port, QN => n_2059
               );
   REGISTERS_reg_31_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N257, 
               clocked_on => CLK_port, Q => REGISTERS_31_17_port, QN => n_2060
               );
   REGISTERS_reg_31_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N256, 
               clocked_on => CLK_port, Q => REGISTERS_31_16_port, QN => n_2061
               );
   REGISTERS_reg_31_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N255, 
               clocked_on => CLK_port, Q => REGISTERS_31_15_port, QN => n_2062
               );
   REGISTERS_reg_31_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N254, 
               clocked_on => CLK_port, Q => REGISTERS_31_14_port, QN => n_2063
               );
   REGISTERS_reg_31_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N253, 
               clocked_on => CLK_port, Q => REGISTERS_31_13_port, QN => n_2064
               );
   REGISTERS_reg_31_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N252, 
               clocked_on => CLK_port, Q => REGISTERS_31_12_port, QN => n_2065
               );
   REGISTERS_reg_31_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N251, 
               clocked_on => CLK_port, Q => REGISTERS_31_11_port, QN => n_2066
               );
   REGISTERS_reg_31_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N250, 
               clocked_on => CLK_port, Q => REGISTERS_31_10_port, QN => n_2067
               );
   REGISTERS_reg_31_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N249, 
               clocked_on => CLK_port, Q => REGISTERS_31_9_port, QN => n_2068);
   REGISTERS_reg_31_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N248, 
               clocked_on => CLK_port, Q => REGISTERS_31_8_port, QN => n_2069);
   REGISTERS_reg_31_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N247, 
               clocked_on => CLK_port, Q => REGISTERS_31_7_port, QN => n_2070);
   REGISTERS_reg_31_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N246, 
               clocked_on => CLK_port, Q => REGISTERS_31_6_port, QN => n_2071);
   REGISTERS_reg_31_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N245, 
               clocked_on => CLK_port, Q => REGISTERS_31_5_port, QN => n_2072);
   REGISTERS_reg_31_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N244, 
               clocked_on => CLK_port, Q => REGISTERS_31_4_port, QN => n_2073);
   REGISTERS_reg_31_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N243, 
               clocked_on => CLK_port, Q => REGISTERS_31_3_port, QN => n_2074);
   REGISTERS_reg_31_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N242, 
               clocked_on => CLK_port, Q => REGISTERS_31_2_port, QN => n_2075);
   REGISTERS_reg_31_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N241, 
               clocked_on => CLK_port, Q => REGISTERS_31_1_port, QN => n_2076);
   REGISTERS_reg_31_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N239, next_state => N240, 
               clocked_on => CLK_port, Q => REGISTERS_31_0_port, QN => n_2077);
   OUT1_reg_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N335, 
               clocked_on => CLK_port, Q => OUT1_31_port, QN => n_2078);
   OUT1_reg_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N334, 
               clocked_on => CLK_port, Q => OUT1_30_port, QN => n_2079);
   OUT1_reg_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N333, 
               clocked_on => CLK_port, Q => OUT1_29_port, QN => n_2080);
   OUT1_reg_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N332, 
               clocked_on => CLK_port, Q => OUT1_28_port, QN => n_2081);
   OUT1_reg_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N331, 
               clocked_on => CLK_port, Q => OUT1_27_port, QN => n_2082);
   OUT1_reg_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N330, 
               clocked_on => CLK_port, Q => OUT1_26_port, QN => n_2083);
   OUT1_reg_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N329, 
               clocked_on => CLK_port, Q => OUT1_25_port, QN => n_2084);
   OUT1_reg_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N328, 
               clocked_on => CLK_port, Q => OUT1_24_port, QN => n_2085);
   OUT1_reg_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N327, 
               clocked_on => CLK_port, Q => OUT1_23_port, QN => n_2086);
   OUT1_reg_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N326, 
               clocked_on => CLK_port, Q => OUT1_22_port, QN => n_2087);
   OUT1_reg_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N325, 
               clocked_on => CLK_port, Q => OUT1_21_port, QN => n_2088);
   OUT1_reg_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N324, 
               clocked_on => CLK_port, Q => OUT1_20_port, QN => n_2089);
   OUT1_reg_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N323, 
               clocked_on => CLK_port, Q => OUT1_19_port, QN => n_2090);
   OUT1_reg_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N322, 
               clocked_on => CLK_port, Q => OUT1_18_port, QN => n_2091);
   OUT1_reg_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N321, 
               clocked_on => CLK_port, Q => OUT1_17_port, QN => n_2092);
   OUT1_reg_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N320, 
               clocked_on => CLK_port, Q => OUT1_16_port, QN => n_2093);
   OUT1_reg_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N319, 
               clocked_on => CLK_port, Q => OUT1_15_port, QN => n_2094);
   OUT1_reg_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N318, 
               clocked_on => CLK_port, Q => OUT1_14_port, QN => n_2095);
   OUT1_reg_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N317, 
               clocked_on => CLK_port, Q => OUT1_13_port, QN => n_2096);
   OUT1_reg_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N316, 
               clocked_on => CLK_port, Q => OUT1_12_port, QN => n_2097);
   OUT1_reg_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N315, 
               clocked_on => CLK_port, Q => OUT1_11_port, QN => n_2098);
   OUT1_reg_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N314, 
               clocked_on => CLK_port, Q => OUT1_10_port, QN => n_2099);
   OUT1_reg_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N313, 
               clocked_on => CLK_port, Q => OUT1_9_port, QN => n_2100);
   OUT1_reg_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N312, 
               clocked_on => CLK_port, Q => OUT1_8_port, QN => n_2101);
   OUT1_reg_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N311, 
               clocked_on => CLK_port, Q => OUT1_7_port, QN => n_2102);
   OUT1_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N310, 
               clocked_on => CLK_port, Q => OUT1_6_port, QN => n_2103);
   OUT1_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N309, 
               clocked_on => CLK_port, Q => OUT1_5_port, QN => n_2104);
   OUT1_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N308, 
               clocked_on => CLK_port, Q => OUT1_4_port, QN => n_2105);
   OUT1_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N307, 
               clocked_on => CLK_port, Q => OUT1_3_port, QN => n_2106);
   OUT1_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N306, 
               clocked_on => CLK_port, Q => OUT1_2_port, QN => n_2107);
   OUT1_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N305, 
               clocked_on => CLK_port, Q => OUT1_1_port, QN => n_2108);
   OUT1_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N303, next_state => N304, 
               clocked_on => CLK_port, Q => OUT1_0_port, QN => n_2109);
   OUT2_reg_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N368, 
               clocked_on => CLK_port, Q => OUT2_31_port, QN => n_2110);
   OUT2_reg_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N367, 
               clocked_on => CLK_port, Q => OUT2_30_port, QN => n_2111);
   OUT2_reg_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N366, 
               clocked_on => CLK_port, Q => OUT2_29_port, QN => n_2112);
   OUT2_reg_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N365, 
               clocked_on => CLK_port, Q => OUT2_28_port, QN => n_2113);
   OUT2_reg_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N364, 
               clocked_on => CLK_port, Q => OUT2_27_port, QN => n_2114);
   OUT2_reg_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N363, 
               clocked_on => CLK_port, Q => OUT2_26_port, QN => n_2115);
   OUT2_reg_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N362, 
               clocked_on => CLK_port, Q => OUT2_25_port, QN => n_2116);
   OUT2_reg_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N361, 
               clocked_on => CLK_port, Q => OUT2_24_port, QN => n_2117);
   OUT2_reg_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N360, 
               clocked_on => CLK_port, Q => OUT2_23_port, QN => n_2118);
   OUT2_reg_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N359, 
               clocked_on => CLK_port, Q => OUT2_22_port, QN => n_2119);
   OUT2_reg_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N358, 
               clocked_on => CLK_port, Q => OUT2_21_port, QN => n_2120);
   OUT2_reg_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N357, 
               clocked_on => CLK_port, Q => OUT2_20_port, QN => n_2121);
   OUT2_reg_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N356, 
               clocked_on => CLK_port, Q => OUT2_19_port, QN => n_2122);
   OUT2_reg_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N355, 
               clocked_on => CLK_port, Q => OUT2_18_port, QN => n_2123);
   OUT2_reg_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N354, 
               clocked_on => CLK_port, Q => OUT2_17_port, QN => n_2124);
   OUT2_reg_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N353, 
               clocked_on => CLK_port, Q => OUT2_16_port, QN => n_2125);
   OUT2_reg_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N352, 
               clocked_on => CLK_port, Q => OUT2_15_port, QN => n_2126);
   OUT2_reg_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N351, 
               clocked_on => CLK_port, Q => OUT2_14_port, QN => n_2127);
   OUT2_reg_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N350, 
               clocked_on => CLK_port, Q => OUT2_13_port, QN => n_2128);
   OUT2_reg_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N349, 
               clocked_on => CLK_port, Q => OUT2_12_port, QN => n_2129);
   OUT2_reg_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N348, 
               clocked_on => CLK_port, Q => OUT2_11_port, QN => n_2130);
   OUT2_reg_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N347, 
               clocked_on => CLK_port, Q => OUT2_10_port, QN => n_2131);
   OUT2_reg_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N346, 
               clocked_on => CLK_port, Q => OUT2_9_port, QN => n_2132);
   OUT2_reg_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N345, 
               clocked_on => CLK_port, Q => OUT2_8_port, QN => n_2133);
   OUT2_reg_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N344, 
               clocked_on => CLK_port, Q => OUT2_7_port, QN => n_2134);
   OUT2_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N343, 
               clocked_on => CLK_port, Q => OUT2_6_port, QN => n_2135);
   OUT2_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N342, 
               clocked_on => CLK_port, Q => OUT2_5_port, QN => n_2136);
   OUT2_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N341, 
               clocked_on => CLK_port, Q => OUT2_4_port, QN => n_2137);
   OUT2_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N340, 
               clocked_on => CLK_port, Q => OUT2_3_port, QN => n_2138);
   OUT2_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N339, 
               clocked_on => CLK_port, Q => OUT2_2_port, QN => n_2139);
   OUT2_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N338, 
               clocked_on => CLK_port, Q => OUT2_1_port, QN => n_2140);
   OUT2_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N336, next_state => N337, 
               clocked_on => CLK_port, Q => OUT2_0_port, QN => n_2141);
   I_0 : GTECH_NOT port map( A => RST, Z => N369);
   C6812 : GTECH_AND2 port map( A => ADD_WR(3), B => ADD_WR(4), Z => N370);
   C6813 : GTECH_AND2 port map( A => N0, B => ADD_WR(4), Z => N371);
   I_1 : GTECH_NOT port map( A => ADD_WR(3), Z => N0);
   C6814 : GTECH_AND2 port map( A => ADD_WR(3), B => N1, Z => N372);
   I_2 : GTECH_NOT port map( A => ADD_WR(4), Z => N1);
   C6815 : GTECH_AND2 port map( A => N2, B => N3, Z => N373);
   I_3 : GTECH_NOT port map( A => ADD_WR(3), Z => N2);
   I_4 : GTECH_NOT port map( A => ADD_WR(4), Z => N3);
   I_5 : GTECH_NOT port map( A => ADD_WR(2), Z => N374);
   C6817 : GTECH_AND2 port map( A => ADD_WR(0), B => ADD_WR(1), Z => N375);
   C6818 : GTECH_AND2 port map( A => N4, B => ADD_WR(1), Z => N376);
   I_6 : GTECH_NOT port map( A => ADD_WR(0), Z => N4);
   C6819 : GTECH_AND2 port map( A => ADD_WR(0), B => N5, Z => N377);
   I_7 : GTECH_NOT port map( A => ADD_WR(1), Z => N5);
   C6820 : GTECH_AND2 port map( A => N6, B => N7, Z => N378);
   I_8 : GTECH_NOT port map( A => ADD_WR(0), Z => N6);
   I_9 : GTECH_NOT port map( A => ADD_WR(1), Z => N7);
   C6821 : GTECH_AND2 port map( A => ADD_WR(2), B => N375, Z => N379);
   C6822 : GTECH_AND2 port map( A => ADD_WR(2), B => N376, Z => N380);
   C6823 : GTECH_AND2 port map( A => ADD_WR(2), B => N377, Z => N381);
   C6824 : GTECH_AND2 port map( A => ADD_WR(2), B => N378, Z => N382);
   C6825 : GTECH_AND2 port map( A => N374, B => N375, Z => N383);
   C6826 : GTECH_AND2 port map( A => N374, B => N376, Z => N384);
   C6827 : GTECH_AND2 port map( A => N374, B => N377, Z => N385);
   C6828 : GTECH_AND2 port map( A => N374, B => N378, Z => N386);
   C6829 : GTECH_AND2 port map( A => N370, B => N379, Z => N387);
   C6830 : GTECH_AND2 port map( A => N370, B => N380, Z => N388);
   C6831 : GTECH_AND2 port map( A => N370, B => N381, Z => N389);
   C6832 : GTECH_AND2 port map( A => N370, B => N382, Z => N390);
   C6833 : GTECH_AND2 port map( A => N370, B => N383, Z => N391);
   C6834 : GTECH_AND2 port map( A => N370, B => N384, Z => N392);
   C6835 : GTECH_AND2 port map( A => N370, B => N385, Z => N393);
   C6836 : GTECH_AND2 port map( A => N370, B => N386, Z => N394);
   C6837 : GTECH_AND2 port map( A => N371, B => N379, Z => N395);
   C6838 : GTECH_AND2 port map( A => N371, B => N380, Z => N396);
   C6839 : GTECH_AND2 port map( A => N371, B => N381, Z => N397);
   C6840 : GTECH_AND2 port map( A => N371, B => N382, Z => N398);
   C6841 : GTECH_AND2 port map( A => N371, B => N383, Z => N399);
   C6842 : GTECH_AND2 port map( A => N371, B => N384, Z => N400);
   C6843 : GTECH_AND2 port map( A => N371, B => N385, Z => N401);
   C6844 : GTECH_AND2 port map( A => N371, B => N386, Z => N402);
   C6845 : GTECH_AND2 port map( A => N372, B => N379, Z => N403);
   C6846 : GTECH_AND2 port map( A => N372, B => N380, Z => N404);
   C6847 : GTECH_AND2 port map( A => N372, B => N381, Z => N405);
   C6848 : GTECH_AND2 port map( A => N372, B => N382, Z => N406);
   C6849 : GTECH_AND2 port map( A => N372, B => N383, Z => N407);
   C6850 : GTECH_AND2 port map( A => N372, B => N384, Z => N408);
   C6851 : GTECH_AND2 port map( A => N372, B => N385, Z => N409);
   C6852 : GTECH_AND2 port map( A => N372, B => N386, Z => N410);
   C6853 : GTECH_AND2 port map( A => N373, B => N379, Z => N411);
   C6854 : GTECH_AND2 port map( A => N373, B => N380, Z => N412);
   C6855 : GTECH_AND2 port map( A => N373, B => N381, Z => N413);
   C6856 : GTECH_AND2 port map( A => N373, B => N382, Z => N414);
   C6857 : GTECH_AND2 port map( A => N373, B => N383, Z => N415);
   C6858 : GTECH_AND2 port map( A => N373, B => N384, Z => N416);
   C6859 : GTECH_AND2 port map( A => N373, B => N385, Z => N417);
   C6860 : GTECH_AND2 port map( A => N373, B => N386, Z => N418);
   C6861_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => N418, DATA(30) => N417, DATA(29) => N416, DATA(28) => N415
               , DATA(27) => N414, DATA(26) => N413, DATA(25) => N412, DATA(24)
               => N411, DATA(23) => N410, DATA(22) => N409, DATA(21) => N408, 
               DATA(20) => N407, DATA(19) => N406, DATA(18) => N405, DATA(17) 
               => N404, DATA(16) => N403, DATA(15) => N402, DATA(14) => N401, 
               DATA(13) => N400, DATA(12) => N399, DATA(11) => N398, DATA(10) 
               => N397, DATA(9) => N396, DATA(8) => N395, DATA(7) => N394, 
               DATA(6) => N393, DATA(5) => N392, DATA(4) => N391, DATA(3) => 
               N390, DATA(2) => N389, DATA(1) => N388, DATA(0) => N387, 
         -- Connections to port 'DATA2'
         DATA(63) => X_Logic0_port, DATA(62) => X_Logic0_port, DATA(61) => 
               X_Logic0_port, DATA(60) => X_Logic0_port, DATA(59) => 
               X_Logic0_port, DATA(58) => X_Logic0_port, DATA(57) => 
               X_Logic0_port, DATA(56) => X_Logic0_port, DATA(55) => 
               X_Logic0_port, DATA(54) => X_Logic0_port, DATA(53) => 
               X_Logic0_port, DATA(52) => X_Logic0_port, DATA(51) => 
               X_Logic0_port, DATA(50) => X_Logic0_port, DATA(49) => 
               X_Logic0_port, DATA(48) => X_Logic0_port, DATA(47) => 
               X_Logic0_port, DATA(46) => X_Logic0_port, DATA(45) => 
               X_Logic0_port, DATA(44) => X_Logic0_port, DATA(43) => 
               X_Logic0_port, DATA(42) => X_Logic0_port, DATA(41) => 
               X_Logic0_port, DATA(40) => X_Logic0_port, DATA(39) => 
               X_Logic0_port, DATA(38) => X_Logic0_port, DATA(37) => 
               X_Logic0_port, DATA(36) => X_Logic0_port, DATA(35) => 
               X_Logic0_port, DATA(34) => X_Logic0_port, DATA(33) => 
               X_Logic0_port, DATA(32) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(31) => N238, Z(30) => N237, Z(29) => N236, Z(28) => N235, Z(27) => 
               N234, Z(26) => N233, Z(25) => N232, Z(24) => N231, Z(23) => N230
               , Z(22) => N229, Z(21) => N228, Z(20) => N227, Z(19) => N226, 
               Z(18) => N225, Z(17) => N224, Z(16) => N223, Z(15) => N222, 
               Z(14) => N221, Z(13) => N220, Z(12) => N219, Z(11) => N218, 
               Z(10) => N217, Z(9) => N216, Z(8) => N215, Z(7) => N214, Z(6) =>
               N213, Z(5) => N212, Z(4) => N211, Z(3) => N210, Z(2) => N209, 
               Z(1) => N208, Z(0) => N207 );
   B_0 : GTECH_BUF port map( A => WR, Z => N8);
   B_1 : GTECH_BUF port map( A => N206, Z => N9);
   C6862_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => X_Logic1_port, DATA(30) => X_Logic1_port, DATA(29) => 
               X_Logic1_port, DATA(28) => X_Logic1_port, DATA(27) => 
               X_Logic1_port, DATA(26) => X_Logic1_port, DATA(25) => 
               X_Logic1_port, DATA(24) => X_Logic1_port, DATA(23) => 
               X_Logic1_port, DATA(22) => X_Logic1_port, DATA(21) => 
               X_Logic1_port, DATA(20) => X_Logic1_port, DATA(19) => 
               X_Logic1_port, DATA(18) => X_Logic1_port, DATA(17) => 
               X_Logic1_port, DATA(16) => X_Logic1_port, DATA(15) => 
               X_Logic1_port, DATA(14) => X_Logic1_port, DATA(13) => 
               X_Logic1_port, DATA(12) => X_Logic1_port, DATA(11) => 
               X_Logic1_port, DATA(10) => X_Logic1_port, DATA(9) => 
               X_Logic1_port, DATA(8) => X_Logic1_port, DATA(7) => 
               X_Logic1_port, DATA(6) => X_Logic1_port, DATA(5) => 
               X_Logic1_port, DATA(4) => X_Logic1_port, DATA(3) => 
               X_Logic1_port, DATA(2) => X_Logic1_port, DATA(1) => 
               X_Logic1_port, DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(63) => N238, DATA(62) => N237, DATA(61) => N236, DATA(60) => N235
               , DATA(59) => N234, DATA(58) => N233, DATA(57) => N232, DATA(56)
               => N231, DATA(55) => N230, DATA(54) => N229, DATA(53) => N228, 
               DATA(52) => N227, DATA(51) => N226, DATA(50) => N225, DATA(49) 
               => N224, DATA(48) => N223, DATA(47) => N222, DATA(46) => N221, 
               DATA(45) => N220, DATA(44) => N219, DATA(43) => N218, DATA(42) 
               => N217, DATA(41) => N216, DATA(40) => N215, DATA(39) => N214, 
               DATA(38) => N213, DATA(37) => N212, DATA(36) => N211, DATA(35) 
               => N210, DATA(34) => N209, DATA(33) => N208, DATA(32) => N207, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(31) => N302, Z(30) => N301, Z(29) => N300, Z(28) => N299, Z(27) => 
               N298, Z(26) => N297, Z(25) => N296, Z(24) => N295, Z(23) => N294
               , Z(22) => N293, Z(21) => N292, Z(20) => N291, Z(19) => N290, 
               Z(18) => N289, Z(17) => N288, Z(16) => N287, Z(15) => N286, 
               Z(14) => N285, Z(13) => N284, Z(12) => N283, Z(11) => N282, 
               Z(10) => N281, Z(9) => N280, Z(8) => N279, Z(7) => N278, Z(6) =>
               N277, Z(5) => N276, Z(4) => N275, Z(3) => N274, Z(2) => N273, 
               Z(1) => N272, Z(0) => N239 );
   B_2 : GTECH_BUF port map( A => N369, Z => N10);
   B_3 : GTECH_BUF port map( A => RST, Z => N11);
   C6863_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => X_Logic0_port, DATA(30) => X_Logic0_port, DATA(29) => 
               X_Logic0_port, DATA(28) => X_Logic0_port, DATA(27) => 
               X_Logic0_port, DATA(26) => X_Logic0_port, DATA(25) => 
               X_Logic0_port, DATA(24) => X_Logic0_port, DATA(23) => 
               X_Logic0_port, DATA(22) => X_Logic0_port, DATA(21) => 
               X_Logic0_port, DATA(20) => X_Logic0_port, DATA(19) => 
               X_Logic0_port, DATA(18) => X_Logic0_port, DATA(17) => 
               X_Logic0_port, DATA(16) => X_Logic0_port, DATA(15) => 
               X_Logic0_port, DATA(14) => X_Logic0_port, DATA(13) => 
               X_Logic0_port, DATA(12) => X_Logic0_port, DATA(11) => 
               X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic0_port, DATA(8) => X_Logic0_port, DATA(7) => 
               X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => DATAIN_31_port, DATA(62) => DATAIN_30_port, DATA(61) => 
               DATAIN_29_port, DATA(60) => DATAIN_28_port, DATA(59) => 
               DATAIN_27_port, DATA(58) => DATAIN_26_port, DATA(57) => 
               DATAIN_25_port, DATA(56) => DATAIN_24_port, DATA(55) => 
               DATAIN_23_port, DATA(54) => DATAIN_22_port, DATA(53) => 
               DATAIN_21_port, DATA(52) => DATAIN_20_port, DATA(51) => 
               DATAIN_19_port, DATA(50) => DATAIN_18_port, DATA(49) => 
               DATAIN_17_port, DATA(48) => DATAIN_16_port, DATA(47) => 
               DATAIN_15_port, DATA(46) => DATAIN_14_port, DATA(45) => 
               DATAIN_13_port, DATA(44) => DATAIN_12_port, DATA(43) => 
               DATAIN_11_port, DATA(42) => DATAIN_10_port, DATA(41) => 
               DATAIN_9_port, DATA(40) => DATAIN_8_port, DATA(39) => 
               DATAIN_7_port, DATA(38) => DATAIN_6_port, DATA(37) => 
               DATAIN_5_port, DATA(36) => DATAIN_4_port, DATA(35) => 
               DATAIN_3_port, DATA(34) => DATAIN_2_port, DATA(33) => 
               DATAIN_1_port, DATA(32) => DATAIN_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(31) => N271, Z(30) => N270, Z(29) => N269, Z(28) => N268, Z(27) => 
               N267, Z(26) => N266, Z(25) => N265, Z(24) => N264, Z(23) => N263
               , Z(22) => N262, Z(21) => N261, Z(20) => N260, Z(19) => N259, 
               Z(18) => N258, Z(17) => N257, Z(16) => N256, Z(15) => N255, 
               Z(14) => N254, Z(13) => N253, Z(12) => N252, Z(11) => N251, 
               Z(10) => N250, Z(9) => N249, Z(8) => N248, Z(7) => N247, Z(6) =>
               N246, Z(5) => N245, Z(4) => N244, Z(3) => N243, Z(2) => N242, 
               Z(1) => N241, Z(0) => N240 );
   C6864_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => RD1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(0) => N303 );
   C6865_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => X_Logic0_port, DATA(30) => X_Logic0_port, DATA(29) => 
               X_Logic0_port, DATA(28) => X_Logic0_port, DATA(27) => 
               X_Logic0_port, DATA(26) => X_Logic0_port, DATA(25) => 
               X_Logic0_port, DATA(24) => X_Logic0_port, DATA(23) => 
               X_Logic0_port, DATA(22) => X_Logic0_port, DATA(21) => 
               X_Logic0_port, DATA(20) => X_Logic0_port, DATA(19) => 
               X_Logic0_port, DATA(18) => X_Logic0_port, DATA(17) => 
               X_Logic0_port, DATA(16) => X_Logic0_port, DATA(15) => 
               X_Logic0_port, DATA(14) => X_Logic0_port, DATA(13) => 
               X_Logic0_port, DATA(12) => X_Logic0_port, DATA(11) => 
               X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic0_port, DATA(8) => X_Logic0_port, DATA(7) => 
               X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => N77, DATA(62) => N78, DATA(61) => N79, DATA(60) => N80, 
               DATA(59) => N81, DATA(58) => N82, DATA(57) => N83, DATA(56) => 
               N84, DATA(55) => N85, DATA(54) => N86, DATA(53) => N87, DATA(52)
               => N88, DATA(51) => N89, DATA(50) => N90, DATA(49) => N91, 
               DATA(48) => N92, DATA(47) => N93, DATA(46) => N94, DATA(45) => 
               N95, DATA(44) => N96, DATA(43) => N97, DATA(42) => N98, DATA(41)
               => N99, DATA(40) => N100, DATA(39) => N101, DATA(38) => N102, 
               DATA(37) => N103, DATA(36) => N104, DATA(35) => N105, DATA(34) 
               => N106, DATA(33) => N107, DATA(32) => N108, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(31) => N335, Z(30) => N334, Z(29) => N333, Z(28) => N332, Z(27) => 
               N331, Z(26) => N330, Z(25) => N329, Z(24) => N328, Z(23) => N327
               , Z(22) => N326, Z(21) => N325, Z(20) => N324, Z(19) => N323, 
               Z(18) => N322, Z(17) => N321, Z(16) => N320, Z(15) => N319, 
               Z(14) => N318, Z(13) => N317, Z(12) => N316, Z(11) => N315, 
               Z(10) => N314, Z(9) => N313, Z(8) => N312, Z(7) => N311, Z(6) =>
               N310, Z(5) => N309, Z(4) => N308, Z(3) => N307, Z(2) => N306, 
               Z(1) => N305, Z(0) => N304 );
   C6866_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => RD2_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(0) => N336 );
   C6867_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => X_Logic0_port, DATA(30) => X_Logic0_port, DATA(29) => 
               X_Logic0_port, DATA(28) => X_Logic0_port, DATA(27) => 
               X_Logic0_port, DATA(26) => X_Logic0_port, DATA(25) => 
               X_Logic0_port, DATA(24) => X_Logic0_port, DATA(23) => 
               X_Logic0_port, DATA(22) => X_Logic0_port, DATA(21) => 
               X_Logic0_port, DATA(20) => X_Logic0_port, DATA(19) => 
               X_Logic0_port, DATA(18) => X_Logic0_port, DATA(17) => 
               X_Logic0_port, DATA(16) => X_Logic0_port, DATA(15) => 
               X_Logic0_port, DATA(14) => X_Logic0_port, DATA(13) => 
               X_Logic0_port, DATA(12) => X_Logic0_port, DATA(11) => 
               X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic0_port, DATA(8) => X_Logic0_port, DATA(7) => 
               X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => N174, DATA(62) => N175, DATA(61) => N176, DATA(60) => N177
               , DATA(59) => N178, DATA(58) => N179, DATA(57) => N180, DATA(56)
               => N181, DATA(55) => N182, DATA(54) => N183, DATA(53) => N184, 
               DATA(52) => N185, DATA(51) => N186, DATA(50) => N187, DATA(49) 
               => N188, DATA(48) => N189, DATA(47) => N190, DATA(46) => N191, 
               DATA(45) => N192, DATA(44) => N193, DATA(43) => N194, DATA(42) 
               => N195, DATA(41) => N196, DATA(40) => N197, DATA(39) => N198, 
               DATA(38) => N199, DATA(37) => N200, DATA(36) => N201, DATA(35) 
               => N202, DATA(34) => N203, DATA(33) => N204, DATA(32) => N205, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(31) => N368, Z(30) => N367, Z(29) => N366, Z(28) => N365, Z(27) => 
               N364, Z(26) => N363, Z(25) => N362, Z(24) => N361, Z(23) => N360
               , Z(22) => N359, Z(21) => N358, Z(20) => N357, Z(19) => N356, 
               Z(18) => N355, Z(17) => N354, Z(16) => N353, Z(15) => N352, 
               Z(14) => N351, Z(13) => N350, Z(12) => N349, Z(11) => N348, 
               Z(10) => N347, Z(9) => N346, Z(8) => N345, Z(7) => N344, Z(6) =>
               N343, Z(5) => N342, Z(4) => N341, Z(3) => N340, Z(2) => N339, 
               Z(1) => N338, Z(0) => N337 );
         X_Logic1_port <= '1';
         X_Logic0_port <= '0';
   I_10 : GTECH_NOT port map( A => ADD_RD1(0), Z => N12);
   I_11 : GTECH_NOT port map( A => ADD_RD1(1), Z => N13);
   C6875 : GTECH_AND2 port map( A => N12, B => N13, Z => N14);
   C6876 : GTECH_AND2 port map( A => N12, B => ADD_RD1(1), Z => N15);
   C6877 : GTECH_AND2 port map( A => ADD_RD1(0), B => N13, Z => N16);
   C6878 : GTECH_AND2 port map( A => ADD_RD1(0), B => ADD_RD1(1), Z => N17);
   I_12 : GTECH_NOT port map( A => ADD_RD1(2), Z => N18);
   C6880 : GTECH_AND2 port map( A => N14, B => N18, Z => N19);
   C6881 : GTECH_AND2 port map( A => N14, B => ADD_RD1(2), Z => N20);
   C6882 : GTECH_AND2 port map( A => N16, B => N18, Z => N21);
   C6883 : GTECH_AND2 port map( A => N16, B => ADD_RD1(2), Z => N22);
   C6884 : GTECH_AND2 port map( A => N15, B => N18, Z => N23);
   C6885 : GTECH_AND2 port map( A => N15, B => ADD_RD1(2), Z => N24);
   C6886 : GTECH_AND2 port map( A => N17, B => N18, Z => N25);
   C6887 : GTECH_AND2 port map( A => N17, B => ADD_RD1(2), Z => N26);
   I_13 : GTECH_NOT port map( A => ADD_RD1(3), Z => N27);
   C6889 : GTECH_AND2 port map( A => N19, B => N27, Z => N28);
   C6890 : GTECH_AND2 port map( A => N19, B => ADD_RD1(3), Z => N29);
   C6891 : GTECH_AND2 port map( A => N21, B => N27, Z => N30);
   C6892 : GTECH_AND2 port map( A => N21, B => ADD_RD1(3), Z => N31);
   C6893 : GTECH_AND2 port map( A => N23, B => N27, Z => N32);
   C6894 : GTECH_AND2 port map( A => N23, B => ADD_RD1(3), Z => N33);
   C6895 : GTECH_AND2 port map( A => N25, B => N27, Z => N34);
   C6896 : GTECH_AND2 port map( A => N25, B => ADD_RD1(3), Z => N35);
   C6897 : GTECH_AND2 port map( A => N20, B => N27, Z => N36);
   C6898 : GTECH_AND2 port map( A => N20, B => ADD_RD1(3), Z => N37);
   C6899 : GTECH_AND2 port map( A => N22, B => N27, Z => N38);
   C6900 : GTECH_AND2 port map( A => N22, B => ADD_RD1(3), Z => N39);
   C6901 : GTECH_AND2 port map( A => N24, B => N27, Z => N40);
   C6902 : GTECH_AND2 port map( A => N24, B => ADD_RD1(3), Z => N41);
   C6903 : GTECH_AND2 port map( A => N26, B => N27, Z => N42);
   C6904 : GTECH_AND2 port map( A => N26, B => ADD_RD1(3), Z => N43);
   I_14 : GTECH_NOT port map( A => ADD_RD1(4), Z => N44);
   C6906 : GTECH_AND2 port map( A => N28, B => N44, Z => N45);
   C6907 : GTECH_AND2 port map( A => N28, B => ADD_RD1(4), Z => N46);
   C6908 : GTECH_AND2 port map( A => N30, B => N44, Z => N47);
   C6909 : GTECH_AND2 port map( A => N30, B => ADD_RD1(4), Z => N48);
   C6910 : GTECH_AND2 port map( A => N32, B => N44, Z => N49);
   C6911 : GTECH_AND2 port map( A => N32, B => ADD_RD1(4), Z => N50);
   C6912 : GTECH_AND2 port map( A => N34, B => N44, Z => N51);
   C6913 : GTECH_AND2 port map( A => N34, B => ADD_RD1(4), Z => N52);
   C6914 : GTECH_AND2 port map( A => N36, B => N44, Z => N53);
   C6915 : GTECH_AND2 port map( A => N36, B => ADD_RD1(4), Z => N54);
   C6916 : GTECH_AND2 port map( A => N38, B => N44, Z => N55);
   C6917 : GTECH_AND2 port map( A => N38, B => ADD_RD1(4), Z => N56);
   C6918 : GTECH_AND2 port map( A => N40, B => N44, Z => N57);
   C6919 : GTECH_AND2 port map( A => N40, B => ADD_RD1(4), Z => N58);
   C6920 : GTECH_AND2 port map( A => N42, B => N44, Z => N59);
   C6921 : GTECH_AND2 port map( A => N42, B => ADD_RD1(4), Z => N60);
   C6922 : GTECH_AND2 port map( A => N29, B => N44, Z => N61);
   C6923 : GTECH_AND2 port map( A => N29, B => ADD_RD1(4), Z => N62);
   C6924 : GTECH_AND2 port map( A => N31, B => N44, Z => N63);
   C6925 : GTECH_AND2 port map( A => N31, B => ADD_RD1(4), Z => N64);
   C6926 : GTECH_AND2 port map( A => N33, B => N44, Z => N65);
   C6927 : GTECH_AND2 port map( A => N33, B => ADD_RD1(4), Z => N66);
   C6928 : GTECH_AND2 port map( A => N35, B => N44, Z => N67);
   C6929 : GTECH_AND2 port map( A => N35, B => ADD_RD1(4), Z => N68);
   C6930 : GTECH_AND2 port map( A => N37, B => N44, Z => N69);
   C6931 : GTECH_AND2 port map( A => N37, B => ADD_RD1(4), Z => N70);
   C6932 : GTECH_AND2 port map( A => N39, B => N44, Z => N71);
   C6933 : GTECH_AND2 port map( A => N39, B => ADD_RD1(4), Z => N72);
   C6934 : GTECH_AND2 port map( A => N41, B => N44, Z => N73);
   C6935 : GTECH_AND2 port map( A => N41, B => ADD_RD1(4), Z => N74);
   C6936 : GTECH_AND2 port map( A => N43, B => N44, Z => N75);
   C6937 : GTECH_AND2 port map( A => N43, B => ADD_RD1(4), Z => N76);
   I_15 : GTECH_NOT port map( A => ADD_RD2(0), Z => N109);
   I_16 : GTECH_NOT port map( A => ADD_RD2(1), Z => N110);
   C6941 : GTECH_AND2 port map( A => N109, B => N110, Z => N111);
   C6942 : GTECH_AND2 port map( A => N109, B => ADD_RD2(1), Z => N112);
   C6943 : GTECH_AND2 port map( A => ADD_RD2(0), B => N110, Z => N113);
   C6944 : GTECH_AND2 port map( A => ADD_RD2(0), B => ADD_RD2(1), Z => N114);
   I_17 : GTECH_NOT port map( A => ADD_RD2(2), Z => N115);
   C6946 : GTECH_AND2 port map( A => N111, B => N115, Z => N116);
   C6947 : GTECH_AND2 port map( A => N111, B => ADD_RD2(2), Z => N117);
   C6948 : GTECH_AND2 port map( A => N113, B => N115, Z => N118);
   C6949 : GTECH_AND2 port map( A => N113, B => ADD_RD2(2), Z => N119);
   C6950 : GTECH_AND2 port map( A => N112, B => N115, Z => N120);
   C6951 : GTECH_AND2 port map( A => N112, B => ADD_RD2(2), Z => N121);
   C6952 : GTECH_AND2 port map( A => N114, B => N115, Z => N122);
   C6953 : GTECH_AND2 port map( A => N114, B => ADD_RD2(2), Z => N123);
   I_18 : GTECH_NOT port map( A => ADD_RD2(3), Z => N124);
   C6955 : GTECH_AND2 port map( A => N116, B => N124, Z => N125);
   C6956 : GTECH_AND2 port map( A => N116, B => ADD_RD2(3), Z => N126);
   C6957 : GTECH_AND2 port map( A => N118, B => N124, Z => N127);
   C6958 : GTECH_AND2 port map( A => N118, B => ADD_RD2(3), Z => N128);
   C6959 : GTECH_AND2 port map( A => N120, B => N124, Z => N129);
   C6960 : GTECH_AND2 port map( A => N120, B => ADD_RD2(3), Z => N130);
   C6961 : GTECH_AND2 port map( A => N122, B => N124, Z => N131);
   C6962 : GTECH_AND2 port map( A => N122, B => ADD_RD2(3), Z => N132);
   C6963 : GTECH_AND2 port map( A => N117, B => N124, Z => N133);
   C6964 : GTECH_AND2 port map( A => N117, B => ADD_RD2(3), Z => N134);
   C6965 : GTECH_AND2 port map( A => N119, B => N124, Z => N135);
   C6966 : GTECH_AND2 port map( A => N119, B => ADD_RD2(3), Z => N136);
   C6967 : GTECH_AND2 port map( A => N121, B => N124, Z => N137);
   C6968 : GTECH_AND2 port map( A => N121, B => ADD_RD2(3), Z => N138);
   C6969 : GTECH_AND2 port map( A => N123, B => N124, Z => N139);
   C6970 : GTECH_AND2 port map( A => N123, B => ADD_RD2(3), Z => N140);
   I_19 : GTECH_NOT port map( A => ADD_RD2(4), Z => N141);
   C6972 : GTECH_AND2 port map( A => N125, B => N141, Z => N142);
   C6973 : GTECH_AND2 port map( A => N125, B => ADD_RD2(4), Z => N143);
   C6974 : GTECH_AND2 port map( A => N127, B => N141, Z => N144);
   C6975 : GTECH_AND2 port map( A => N127, B => ADD_RD2(4), Z => N145);
   C6976 : GTECH_AND2 port map( A => N129, B => N141, Z => N146);
   C6977 : GTECH_AND2 port map( A => N129, B => ADD_RD2(4), Z => N147);
   C6978 : GTECH_AND2 port map( A => N131, B => N141, Z => N148);
   C6979 : GTECH_AND2 port map( A => N131, B => ADD_RD2(4), Z => N149);
   C6980 : GTECH_AND2 port map( A => N133, B => N141, Z => N150);
   C6981 : GTECH_AND2 port map( A => N133, B => ADD_RD2(4), Z => N151);
   C6982 : GTECH_AND2 port map( A => N135, B => N141, Z => N152);
   C6983 : GTECH_AND2 port map( A => N135, B => ADD_RD2(4), Z => N153);
   C6984 : GTECH_AND2 port map( A => N137, B => N141, Z => N154);
   C6985 : GTECH_AND2 port map( A => N137, B => ADD_RD2(4), Z => N155);
   C6986 : GTECH_AND2 port map( A => N139, B => N141, Z => N156);
   C6987 : GTECH_AND2 port map( A => N139, B => ADD_RD2(4), Z => N157);
   C6988 : GTECH_AND2 port map( A => N126, B => N141, Z => N158);
   C6989 : GTECH_AND2 port map( A => N126, B => ADD_RD2(4), Z => N159);
   C6990 : GTECH_AND2 port map( A => N128, B => N141, Z => N160);
   C6991 : GTECH_AND2 port map( A => N128, B => ADD_RD2(4), Z => N161);
   C6992 : GTECH_AND2 port map( A => N130, B => N141, Z => N162);
   C6993 : GTECH_AND2 port map( A => N130, B => ADD_RD2(4), Z => N163);
   C6994 : GTECH_AND2 port map( A => N132, B => N141, Z => N164);
   C6995 : GTECH_AND2 port map( A => N132, B => ADD_RD2(4), Z => N165);
   C6996 : GTECH_AND2 port map( A => N134, B => N141, Z => N166);
   C6997 : GTECH_AND2 port map( A => N134, B => ADD_RD2(4), Z => N167);
   C6998 : GTECH_AND2 port map( A => N136, B => N141, Z => N168);
   C6999 : GTECH_AND2 port map( A => N136, B => ADD_RD2(4), Z => N169);
   C7000 : GTECH_AND2 port map( A => N138, B => N141, Z => N170);
   C7001 : GTECH_AND2 port map( A => N138, B => ADD_RD2(4), Z => N171);
   C7002 : GTECH_AND2 port map( A => N140, B => N141, Z => N172);
   C7003 : GTECH_AND2 port map( A => N140, B => ADD_RD2(4), Z => N173);
   I_20 : GTECH_NOT port map( A => WR, Z => N206);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_N32 is

   port( CURR_ADDR : in std_logic_vector (31 downto 0);  NEXT_ADDR : out 
         std_logic_vector (31 downto 0));

end ADDER_N32;

architecture SYN_BEHAVIOR of ADDER_N32 is

   component ADDER_N32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n3, n_2142 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '1';
   n3 <= '0';
   add_26 : ADDER_N32_DW01_add_0 port map( A(31) => CURR_ADDR(31), A(30) => 
                           CURR_ADDR(30), A(29) => CURR_ADDR(29), A(28) => 
                           CURR_ADDR(28), A(27) => CURR_ADDR(27), A(26) => 
                           CURR_ADDR(26), A(25) => CURR_ADDR(25), A(24) => 
                           CURR_ADDR(24), A(23) => CURR_ADDR(23), A(22) => 
                           CURR_ADDR(22), A(21) => CURR_ADDR(21), A(20) => 
                           CURR_ADDR(20), A(19) => CURR_ADDR(19), A(18) => 
                           CURR_ADDR(18), A(17) => CURR_ADDR(17), A(16) => 
                           CURR_ADDR(16), A(15) => CURR_ADDR(15), A(14) => 
                           CURR_ADDR(14), A(13) => CURR_ADDR(13), A(12) => 
                           CURR_ADDR(12), A(11) => CURR_ADDR(11), A(10) => 
                           CURR_ADDR(10), A(9) => CURR_ADDR(9), A(8) => 
                           CURR_ADDR(8), A(7) => CURR_ADDR(7), A(6) => 
                           CURR_ADDR(6), A(5) => CURR_ADDR(5), A(4) => 
                           CURR_ADDR(4), A(3) => CURR_ADDR(3), A(2) => 
                           CURR_ADDR(2), A(1) => CURR_ADDR(1), A(0) => 
                           CURR_ADDR(0), B(31) => n1, B(30) => n1, B(29) => n1,
                           B(28) => n1, B(27) => n1, B(26) => n1, B(25) => n1, 
                           B(24) => n1, B(23) => n1, B(22) => n1, B(21) => n1, 
                           B(20) => n1, B(19) => n1, B(18) => n1, B(17) => n1, 
                           B(16) => n1, B(15) => n1, B(14) => n1, B(13) => n1, 
                           B(12) => n1, B(11) => n1, B(10) => n1, B(9) => n1, 
                           B(8) => n1, B(7) => n1, B(6) => n1, B(5) => n1, B(4)
                           => n1, B(3) => n1, B(2) => n2, B(1) => n1, B(0) => 
                           n1, CI => n3, SUM(31) => NEXT_ADDR(31), SUM(30) => 
                           NEXT_ADDR(30), SUM(29) => NEXT_ADDR(29), SUM(28) => 
                           NEXT_ADDR(28), SUM(27) => NEXT_ADDR(27), SUM(26) => 
                           NEXT_ADDR(26), SUM(25) => NEXT_ADDR(25), SUM(24) => 
                           NEXT_ADDR(24), SUM(23) => NEXT_ADDR(23), SUM(22) => 
                           NEXT_ADDR(22), SUM(21) => NEXT_ADDR(21), SUM(20) => 
                           NEXT_ADDR(20), SUM(19) => NEXT_ADDR(19), SUM(18) => 
                           NEXT_ADDR(18), SUM(17) => NEXT_ADDR(17), SUM(16) => 
                           NEXT_ADDR(16), SUM(15) => NEXT_ADDR(15), SUM(14) => 
                           NEXT_ADDR(14), SUM(13) => NEXT_ADDR(13), SUM(12) => 
                           NEXT_ADDR(12), SUM(11) => NEXT_ADDR(11), SUM(10) => 
                           NEXT_ADDR(10), SUM(9) => NEXT_ADDR(9), SUM(8) => 
                           NEXT_ADDR(8), SUM(7) => NEXT_ADDR(7), SUM(6) => 
                           NEXT_ADDR(6), SUM(5) => NEXT_ADDR(5), SUM(4) => 
                           NEXT_ADDR(4), SUM(3) => NEXT_ADDR(3), SUM(2) => 
                           NEXT_ADDR(2), SUM(1) => NEXT_ADDR(1), SUM(0) => 
                           NEXT_ADDR(0), CO => n_2142);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT5_0 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_GENERIC_NBIT5_0;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT5_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U5 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21 is

   port( A, B, SEL : in std_logic;  Y : out std_logic);

end MUX21;

architecture SYN_BEHAVIOR of MUX21 is

   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X2 port map( A => A, B => B, S => SEL, Z => Y);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_0;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BRANCHING_UNIT_N32 is

   port( CLK, RST : in std_logic;  Reg_A : in std_logic_vector (31 downto 0);  
         EQ_cond, IS_JUMP : in std_logic;  branch_taken : out std_logic);

end BRANCHING_UNIT_N32;

architecture SYN_BEHAVIOR of BRANCHING_UNIT_N32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n_2143 :
      std_logic;

begin
   
   branch_taken_reg : DFF_X1 port map( D => n14, CK => CLK, Q => branch_taken, 
                           QN => n_2143);
   U3 : INV_X1 port map( A => n1, ZN => n14);
   U4 : OAI21_X1 port map( B1 => IS_JUMP, B2 => n2, A => RST, ZN => n1);
   U5 : XNOR2_X1 port map( A => EQ_cond, B => n3, ZN => n2);
   U6 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n3);
   U7 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n5);
   U8 : NOR4_X1 port map( A1 => Reg_A(23), A2 => Reg_A(22), A3 => Reg_A(21), A4
                           => Reg_A(20), ZN => n9);
   U9 : NOR4_X1 port map( A1 => Reg_A(1), A2 => Reg_A(19), A3 => Reg_A(18), A4 
                           => Reg_A(17), ZN => n8);
   U10 : NOR4_X1 port map( A1 => Reg_A(16), A2 => Reg_A(15), A3 => Reg_A(14), 
                           A4 => Reg_A(13), ZN => n7);
   U11 : NOR4_X1 port map( A1 => Reg_A(12), A2 => Reg_A(11), A3 => Reg_A(10), 
                           A4 => Reg_A(0), ZN => n6);
   U12 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12, A4 => n13, ZN => 
                           n4);
   U13 : NOR4_X1 port map( A1 => Reg_A(9), A2 => Reg_A(8), A3 => Reg_A(7), A4 
                           => Reg_A(6), ZN => n13);
   U14 : NOR4_X1 port map( A1 => Reg_A(5), A2 => Reg_A(4), A3 => Reg_A(3), A4 
                           => Reg_A(31), ZN => n12);
   U15 : NOR4_X1 port map( A1 => Reg_A(30), A2 => Reg_A(2), A3 => Reg_A(29), A4
                           => Reg_A(28), ZN => n11);
   U16 : NOR4_X1 port map( A1 => Reg_A(27), A2 => Reg_A(26), A3 => Reg_A(25), 
                           A4 => Reg_A(24), ZN => n10);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT5_0 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 downto 
         0);  DATA_OUT : out std_logic_vector (4 downto 0));

end REG_GENERIC_NBIT5_0;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n14, CK => CLK, Q => DATA_OUT(4)
                           , QN => n13);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n15, CK => CLK, Q => DATA_OUT(3)
                           , QN => n12);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n16, CK => CLK, Q => DATA_OUT(2)
                           , QN => n11);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n17, CK => CLK, Q => DATA_OUT(1)
                           , QN => n10);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n18, CK => CLK, Q => DATA_OUT(0)
                           , QN => n9);
   U3 : OAI21_X1 port map( B1 => n13, B2 => n1, A => n2, ZN => n14);
   U4 : NAND2_X1 port map( A1 => DATA_IN(4), A2 => n3, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n12, B2 => n1, A => n4, ZN => n15);
   U6 : NAND2_X1 port map( A1 => DATA_IN(3), A2 => n3, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n11, B2 => n1, A => n5, ZN => n16);
   U8 : NAND2_X1 port map( A1 => DATA_IN(2), A2 => n3, ZN => n5);
   U9 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n6, ZN => n17);
   U10 : NAND2_X1 port map( A1 => DATA_IN(1), A2 => n3, ZN => n6);
   U11 : OAI21_X1 port map( B1 => n9, B2 => n1, A => n7, ZN => n18);
   U12 : NAND2_X1 port map( A1 => DATA_IN(0), A2 => n3, ZN => n7);
   U13 : AND2_X1 port map( A1 => RST, A2 => n1, ZN => n3);
   U14 : NAND2_X1 port map( A1 => n8, A2 => RST, ZN => n1);
   U15 : INV_X1 port map( A => EN, ZN => n8);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT16 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (15 downto
         0);  DATA_OUT : out std_logic_vector (15 downto 0));

end REG_GENERIC_NBIT16;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51 : std_logic;

begin
   
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n36, CK => CLK, Q => 
                           DATA_OUT(15), QN => n35);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n37, CK => CLK, Q => 
                           DATA_OUT(14), QN => n34);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n38, CK => CLK, Q => 
                           DATA_OUT(13), QN => n33);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n39, CK => CLK, Q => 
                           DATA_OUT(12), QN => n32);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n40, CK => CLK, Q => 
                           DATA_OUT(11), QN => n31);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n41, CK => CLK, Q => 
                           DATA_OUT(10), QN => n30);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n42, CK => CLK, Q => DATA_OUT(9)
                           , QN => n29);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n43, CK => CLK, Q => DATA_OUT(8)
                           , QN => n28);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n44, CK => CLK, Q => DATA_OUT(7)
                           , QN => n27);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n45, CK => CLK, Q => DATA_OUT(6)
                           , QN => n26);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n46, CK => CLK, Q => DATA_OUT(5)
                           , QN => n25);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n47, CK => CLK, Q => DATA_OUT(4)
                           , QN => n24);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n48, CK => CLK, Q => DATA_OUT(3)
                           , QN => n23);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n49, CK => CLK, Q => DATA_OUT(2)
                           , QN => n22);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n50, CK => CLK, Q => DATA_OUT(1)
                           , QN => n21);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n51, CK => CLK, Q => DATA_OUT(0)
                           , QN => n20);
   U3 : OAI22_X1 port map( A1 => n35, A2 => n1, B1 => n2, B2 => n3, ZN => n36);
   U4 : INV_X1 port map( A => DATA_IN(15), ZN => n3);
   U5 : OAI22_X1 port map( A1 => n34, A2 => n1, B1 => n2, B2 => n4, ZN => n37);
   U6 : INV_X1 port map( A => DATA_IN(14), ZN => n4);
   U7 : OAI22_X1 port map( A1 => n33, A2 => n1, B1 => n2, B2 => n5, ZN => n38);
   U8 : INV_X1 port map( A => DATA_IN(13), ZN => n5);
   U9 : OAI22_X1 port map( A1 => n32, A2 => n1, B1 => n2, B2 => n6, ZN => n39);
   U10 : INV_X1 port map( A => DATA_IN(12), ZN => n6);
   U11 : OAI22_X1 port map( A1 => n31, A2 => n1, B1 => n2, B2 => n7, ZN => n40)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(11), ZN => n7);
   U13 : OAI22_X1 port map( A1 => n30, A2 => n1, B1 => n2, B2 => n8, ZN => n41)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(10), ZN => n8);
   U15 : OAI22_X1 port map( A1 => n29, A2 => n1, B1 => n2, B2 => n9, ZN => n42)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(9), ZN => n9);
   U17 : OAI22_X1 port map( A1 => n28, A2 => n1, B1 => n2, B2 => n10, ZN => n43
                           );
   U18 : INV_X1 port map( A => DATA_IN(8), ZN => n10);
   U19 : OAI22_X1 port map( A1 => n27, A2 => n1, B1 => n2, B2 => n11, ZN => n44
                           );
   U20 : INV_X1 port map( A => DATA_IN(7), ZN => n11);
   U21 : OAI22_X1 port map( A1 => n26, A2 => n1, B1 => n2, B2 => n12, ZN => n45
                           );
   U22 : INV_X1 port map( A => DATA_IN(6), ZN => n12);
   U23 : OAI22_X1 port map( A1 => n25, A2 => n1, B1 => n2, B2 => n13, ZN => n46
                           );
   U24 : INV_X1 port map( A => DATA_IN(5), ZN => n13);
   U25 : OAI22_X1 port map( A1 => n24, A2 => n1, B1 => n2, B2 => n14, ZN => n47
                           );
   U26 : INV_X1 port map( A => DATA_IN(4), ZN => n14);
   U27 : OAI22_X1 port map( A1 => n23, A2 => n1, B1 => n2, B2 => n15, ZN => n48
                           );
   U28 : INV_X1 port map( A => DATA_IN(3), ZN => n15);
   U29 : OAI22_X1 port map( A1 => n22, A2 => n1, B1 => n2, B2 => n16, ZN => n49
                           );
   U30 : INV_X1 port map( A => DATA_IN(2), ZN => n16);
   U31 : OAI22_X1 port map( A1 => n21, A2 => n1, B1 => n2, B2 => n17, ZN => n50
                           );
   U32 : INV_X1 port map( A => DATA_IN(1), ZN => n17);
   U33 : OAI22_X1 port map( A1 => n20, A2 => n1, B1 => n2, B2 => n18, ZN => n51
                           );
   U34 : INV_X1 port map( A => DATA_IN(0), ZN => n18);
   U35 : NAND2_X1 port map( A1 => RST, A2 => n1, ZN => n2);
   U36 : NAND2_X1 port map( A1 => n19, A2 => RST, ZN => n1);
   U37 : INV_X1 port map( A => EN, ZN => n19);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity dlx_cu is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
         EQ_COND, IS_JUMP : out std_logic;  ALU_OPCODE : out std_logic_vector 
         (0 to 3);  DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, IS_JAL, 
         WB_MUX_SEL, RF_WE : out std_logic);

end dlx_cu;

architecture SYN_dlx_cu_hw of dlx_cu is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal aluOpcode1_3_port, aluOpcode1_2_port, aluOpcode1_1_port, 
      aluOpcode1_0_port, aluOpcode_i_3_port, aluOpcode_i_2_port, 
      aluOpcode_i_1_port, aluOpcode_i_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, 
      n_2150, n_2151 : std_logic;

begin
   
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_3_port, QN => n_2144);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_2_port, QN => n_2145);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_1_port, QN => n_2146);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_0_port, QN => n_2147);
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => aluOpcode1_3_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(0), QN => n_2148);
   aluOpcode2_reg_2_inst : DFFR_X1 port map( D => aluOpcode1_2_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(1), QN => n_2149);
   aluOpcode2_reg_1_inst : DFFR_X1 port map( D => aluOpcode1_1_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(2), QN => n_2150);
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => aluOpcode1_0_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(3), QN => n_2151);
   RF_WE <= '0';
   WB_MUX_SEL <= '0';
   IS_JAL <= '0';
   PC_LATCH_EN <= '0';
   JUMP_EN <= '0';
   LMD_LATCH_EN <= '0';
   DRAM_WE <= '0';
   IS_JUMP <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   NPC_LATCH_EN <= '0';
   IR_LATCH_EN <= '0';
   SIGNED_IMM <= '0';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   U21 : OAI211_X1 port map( C1 => n1, C2 => n2, A => n3, B => n4, ZN => 
                           aluOpcode_i_3_port);
   U22 : INV_X1 port map( A => n5, ZN => n4);
   U23 : OAI22_X1 port map( A1 => n6, A2 => IR_IN(2), B1 => n7, B2 => IR_IN(28)
                           , ZN => n5);
   U24 : INV_X1 port map( A => n8, ZN => n2);
   U25 : OAI211_X1 port map( C1 => n9, C2 => n10, A => n11, B => n12, ZN => 
                           aluOpcode_i_2_port);
   U26 : NAND4_X1 port map( A1 => n13, A2 => n14, A3 => IR_IN(2), A4 => n15, ZN
                           => n11);
   U27 : INV_X1 port map( A => n16, ZN => n15);
   U28 : XNOR2_X1 port map( A => IR_IN(1), B => n17, ZN => n13);
   U29 : NOR2_X1 port map( A1 => IR_IN(0), A2 => IR_IN(3), ZN => n17);
   U30 : MUX2_X1 port map( A => n18, B => n19, S => n20, Z => n10);
   U31 : AOI22_X1 port map( A1 => n21, A2 => IR_IN(28), B1 => IR_IN(27), B2 => 
                           n22, ZN => n19);
   U32 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => n18);
   U33 : INV_X1 port map( A => n24, ZN => aluOpcode_i_1_port);
   U34 : AOI211_X1 port map( C1 => n8, C2 => n25, A => n26, B => n27, ZN => n24
                           );
   U35 : OAI33_X1 port map( A1 => n28, A2 => IR_IN(27), A3 => n29, B1 => n30, 
                           B2 => n9, B3 => n31, ZN => n26);
   U36 : INV_X1 port map( A => n32, ZN => n31);
   U37 : OR3_X1 port map( A1 => IR_IN(30), A2 => IR_IN(31), A3 => IR_IN(26), ZN
                           => n30);
   U38 : OAI21_X1 port map( B1 => IR_IN(1), B2 => n33, A => n34, ZN => n25);
   U39 : NAND3_X1 port map( A1 => n14, A2 => n35, A3 => n36, ZN => n34);
   U40 : INV_X1 port map( A => IR_IN(3), ZN => n35);
   U41 : AOI21_X1 port map( B1 => n14, B2 => IR_IN(2), A => n37, ZN => n33);
   U42 : INV_X1 port map( A => n38, ZN => n14);
   U43 : OAI211_X1 port map( C1 => n23, C2 => n3, A => n12, B => n39, ZN => 
                           aluOpcode_i_0_port);
   U44 : AOI22_X1 port map( A1 => n8, A2 => n40, B1 => n41, B2 => n20, ZN => 
                           n39);
   U45 : INV_X1 port map( A => IR_IN(30), ZN => n20);
   U46 : OAI21_X1 port map( B1 => n28, B2 => n9, A => n42, ZN => n41);
   U47 : MUX2_X1 port map( A => n43, B => n44, S => IR_IN(31), Z => n42);
   U48 : NAND2_X1 port map( A1 => n32, A2 => IR_IN(26), ZN => n44);
   U49 : MUX2_X1 port map( A => n45, B => n46, S => n9, Z => n43);
   U50 : AOI21_X1 port map( B1 => IR_IN(28), B2 => n23, A => n32, ZN => n46);
   U51 : NOR2_X1 port map( A1 => n23, A2 => IR_IN(28), ZN => n32);
   U52 : NAND2_X1 port map( A1 => n47, A2 => n23, ZN => n45);
   U53 : INV_X1 port map( A => n22, ZN => n28);
   U54 : OAI22_X1 port map( A1 => n1, A2 => n48, B1 => n38, B2 => n49, ZN => 
                           n40);
   U55 : OR2_X1 port map( A1 => n36, A2 => IR_IN(3), ZN => n49);
   U56 : NOR2_X1 port map( A1 => n48, A2 => IR_IN(2), ZN => n36);
   U57 : INV_X1 port map( A => IR_IN(1), ZN => n48);
   U58 : INV_X1 port map( A => n37, ZN => n1);
   U59 : NOR4_X1 port map( A1 => n50, A2 => n51, A3 => IR_IN(3), A4 => IR_IN(5)
                           , ZN => n37);
   U60 : INV_X1 port map( A => n52, ZN => n51);
   U61 : NOR2_X1 port map( A1 => n16, A2 => IR_IN(0), ZN => n8);
   U62 : INV_X1 port map( A => n27, ZN => n12);
   U63 : OAI22_X1 port map( A1 => n53, A2 => n7, B1 => n50, B2 => n6, ZN => n27
                           );
   U64 : NAND3_X1 port map( A1 => IR_IN(3), A2 => IR_IN(0), A3 => n54, ZN => n6
                           );
   U65 : NOR3_X1 port map( A1 => n38, A2 => IR_IN(1), A3 => n16, ZN => n54);
   U66 : NAND4_X1 port map( A1 => n29, A2 => n47, A3 => n55, A4 => n23, ZN => 
                           n16);
   U67 : NOR2_X1 port map( A1 => IR_IN(31), A2 => IR_IN(28), ZN => n55);
   U68 : NOR2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), ZN => n29);
   U69 : NAND2_X1 port map( A1 => IR_IN(5), A2 => n52, ZN => n38);
   U70 : NOR4_X1 port map( A1 => IR_IN(6), A2 => IR_IN(4), A3 => IR_IN(10), A4 
                           => n56, ZN => n52);
   U71 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN =>
                           n56);
   U72 : INV_X1 port map( A => IR_IN(2), ZN => n50);
   U73 : NAND3_X1 port map( A1 => n21, A2 => IR_IN(30), A3 => IR_IN(29), ZN => 
                           n7);
   U74 : NOR3_X1 port map( A1 => IR_IN(27), A2 => IR_IN(31), A3 => n47, ZN => 
                           n21);
   U75 : INV_X1 port map( A => IR_IN(26), ZN => n47);
   U76 : NAND3_X1 port map( A1 => n22, A2 => n9, A3 => IR_IN(30), ZN => n3);
   U77 : INV_X1 port map( A => IR_IN(29), ZN => n9);
   U78 : NOR3_X1 port map( A1 => IR_IN(26), A2 => IR_IN(31), A3 => n53, ZN => 
                           n22);
   U79 : INV_X1 port map( A => IR_IN(28), ZN => n53);
   U80 : INV_X1 port map( A => IR_IN(27), ZN => n23);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 is

   port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
         EQ_COND, IS_JUMP : in std_logic;  ALU_OPCODE : in std_logic_vector (0 
         to 3);  JUMP_EN, PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE : in std_logic
         ;  D_ADDR : out std_logic_vector (5 downto 0);  D_DATA_IN : out 
         std_logic_vector (31 downto 0);  D_DATA_OUT, PC_IN : in 
         std_logic_vector (31 downto 0);  PC_BUS : out std_logic_vector (31 
         downto 0));

end DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64;

architecture SYN_STRUCTURE of 
   DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component ALU_N32
      port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component EXTENDER_NBIT32_IMM_field_lenght16
      port( NOT_EXT_IMM : in std_logic_vector (15 downto 0);  SIGNED_IMM : in 
            std_logic;  EXT_IMM : out std_logic_vector (31 downto 0));
   end component;
   
   component ADDER_N32
      port( CURR_ADDR : in std_logic_vector (31 downto 0);  NEXT_ADDR : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT5_1
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT5_0
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component MUX21
      port( A, B, SEL : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component BRANCHING_UNIT_N32
      port( CLK, RST : in std_logic;  Reg_A : in std_logic_vector (31 downto 0)
            ;  EQ_cond, IS_JUMP : in std_logic;  branch_taken : out std_logic);
   end component;
   
   component REG_GENERIC_NBIT32_1
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_2
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_3
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT5_1
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 
            downto 0);  DATA_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component REG_GENERIC_NBIT5_2
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 
            downto 0);  DATA_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component REG_GENERIC_NBIT5_0
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 
            downto 0);  DATA_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component REG_GENERIC_NBIT16
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (15 
            downto 0);  DATA_OUT : out std_logic_vector (15 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_4
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_5
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_6
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_7
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_8
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REGISTER_FILE_NBIT32_NREG32
      port( CLK, RST, EN, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, D_ADDR_5_port, D_ADDR_4_port, 
      D_ADDR_3_port, D_ADDR_2_port, D_ADDR_1_port, D_ADDR_0_port, 
      PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, current_PC_31_port, 
      current_PC_30_port, current_PC_29_port, current_PC_28_port, 
      current_PC_27_port, current_PC_26_port, current_PC_25_port, 
      current_PC_24_port, current_PC_23_port, current_PC_22_port, 
      current_PC_21_port, current_PC_20_port, current_PC_19_port, 
      current_PC_18_port, current_PC_17_port, current_PC_16_port, 
      current_PC_15_port, current_PC_14_port, current_PC_13_port, 
      current_PC_12_port, current_PC_11_port, current_PC_10_port, 
      current_PC_9_port, current_PC_8_port, current_PC_7_port, 
      current_PC_6_port, current_PC_5_port, current_PC_4_port, 
      current_PC_3_port, current_PC_2_port, current_PC_1_port, 
      current_PC_0_port, current_PC1_31_port, current_PC1_30_port, 
      current_PC1_29_port, current_PC1_28_port, current_PC1_27_port, 
      current_PC1_26_port, current_PC1_25_port, current_PC1_24_port, 
      current_PC1_23_port, current_PC1_22_port, current_PC1_21_port, 
      current_PC1_20_port, current_PC1_19_port, current_PC1_18_port, 
      current_PC1_17_port, current_PC1_16_port, current_PC1_15_port, 
      current_PC1_14_port, current_PC1_13_port, current_PC1_12_port, 
      current_PC1_11_port, current_PC1_10_port, current_PC1_9_port, 
      current_PC1_8_port, current_PC1_7_port, current_PC1_6_port, 
      current_PC1_5_port, current_PC1_4_port, current_PC1_3_port, 
      current_PC1_2_port, current_PC1_1_port, current_PC1_0_port, 
      current_PC2_31_port, current_PC2_30_port, current_PC2_29_port, 
      current_PC2_28_port, current_PC2_27_port, current_PC2_26_port, 
      current_PC2_25_port, current_PC2_24_port, current_PC2_23_port, 
      current_PC2_22_port, current_PC2_21_port, current_PC2_20_port, 
      current_PC2_19_port, current_PC2_18_port, current_PC2_17_port, 
      current_PC2_16_port, current_PC2_15_port, current_PC2_14_port, 
      current_PC2_13_port, current_PC2_12_port, current_PC2_11_port, 
      current_PC2_10_port, current_PC2_9_port, current_PC2_8_port, 
      current_PC2_7_port, current_PC2_6_port, current_PC2_5_port, 
      current_PC2_4_port, current_PC2_3_port, current_PC2_2_port, 
      current_PC2_1_port, current_PC2_0_port, current_PC3_31_port, 
      current_PC3_30_port, current_PC3_29_port, current_PC3_28_port, 
      current_PC3_27_port, current_PC3_26_port, current_PC3_25_port, 
      current_PC3_24_port, current_PC3_23_port, current_PC3_22_port, 
      current_PC3_21_port, current_PC3_20_port, current_PC3_19_port, 
      current_PC3_18_port, current_PC3_17_port, current_PC3_16_port, 
      current_PC3_15_port, current_PC3_14_port, current_PC3_13_port, 
      current_PC3_12_port, current_PC3_11_port, current_PC3_10_port, 
      current_PC3_9_port, current_PC3_8_port, current_PC3_7_port, 
      current_PC3_6_port, current_PC3_5_port, current_PC3_4_port, 
      current_PC3_3_port, current_PC3_2_port, current_PC3_1_port, 
      current_PC3_0_port, next_NPC_31_port, next_NPC_30_port, next_NPC_29_port,
      next_NPC_28_port, next_NPC_27_port, next_NPC_26_port, next_NPC_25_port, 
      next_NPC_24_port, next_NPC_23_port, next_NPC_22_port, next_NPC_21_port, 
      next_NPC_20_port, next_NPC_19_port, next_NPC_18_port, next_NPC_17_port, 
      next_NPC_16_port, next_NPC_15_port, next_NPC_14_port, next_NPC_13_port, 
      next_NPC_12_port, next_NPC_11_port, next_NPC_10_port, next_NPC_9_port, 
      next_NPC_8_port, next_NPC_7_port, next_NPC_6_port, next_NPC_5_port, 
      next_NPC_4_port, next_NPC_3_port, next_NPC_2_port, next_NPC_1_port, 
      next_NPC_0_port, current_NPC_31_port, current_NPC_30_port, 
      current_NPC_29_port, current_NPC_28_port, current_NPC_27_port, 
      current_NPC_26_port, current_NPC_25_port, current_NPC_24_port, 
      current_NPC_23_port, current_NPC_22_port, current_NPC_21_port, 
      current_NPC_20_port, current_NPC_19_port, current_NPC_18_port, 
      current_NPC_17_port, current_NPC_16_port, current_NPC_15_port, 
      current_NPC_14_port, current_NPC_13_port, current_NPC_12_port, 
      current_NPC_11_port, current_NPC_10_port, current_NPC_9_port, 
      current_NPC_8_port, current_NPC_7_port, current_NPC_6_port, 
      current_NPC_5_port, current_NPC_4_port, current_NPC_3_port, 
      current_NPC_2_port, current_NPC_1_port, current_NPC_0_port, 
      current_IW_25_port, current_IW_24_port, current_IW_23_port, 
      current_IW_22_port, current_IW_21_port, current_IW_20_port, 
      current_IW_19_port, current_IW_18_port, current_IW_17_port, 
      current_IW_16_port, current_IW_15_port, current_IW_14_port, 
      current_IW_13_port, current_IW_12_port, current_IW_11_port, 
      current_IW_10_port, current_IW_9_port, current_IW_8_port, 
      current_IW_7_port, current_IW_6_port, current_IW_5_port, 
      current_IW_4_port, current_IW_3_port, current_IW_2_port, 
      current_IW_1_port, current_IW_0_port, IMM_IN_15_port, IMM_IN_14_port, 
      IMM_IN_13_port, IMM_IN_12_port, IMM_IN_11_port, IMM_IN_10_port, 
      IMM_IN_9_port, IMM_IN_8_port, IMM_IN_7_port, IMM_IN_6_port, IMM_IN_5_port
      , IMM_IN_4_port, IMM_IN_3_port, IMM_IN_2_port, IMM_IN_1_port, 
      IMM_IN_0_port, WB1_IN_4_port, WB1_IN_3_port, WB1_IN_2_port, WB1_IN_1_port
      , WB1_IN_0_port, WB2_IN_4_port, WB2_IN_3_port, WB2_IN_2_port, 
      WB2_IN_1_port, WB2_IN_0_port, WB2_OUT_4_port, WB2_OUT_3_port, 
      WB2_OUT_2_port, WB2_OUT_1_port, WB2_OUT_0_port, WB3_OUT_4_port, 
      WB3_OUT_3_port, WB3_OUT_2_port, WB3_OUT_1_port, WB3_OUT_0_port, 
      next_ALU_OUT_31_port, next_ALU_OUT_30_port, next_ALU_OUT_29_port, 
      next_ALU_OUT_28_port, next_ALU_OUT_27_port, next_ALU_OUT_26_port, 
      next_ALU_OUT_25_port, next_ALU_OUT_24_port, next_ALU_OUT_23_port, 
      next_ALU_OUT_22_port, next_ALU_OUT_21_port, next_ALU_OUT_20_port, 
      next_ALU_OUT_19_port, next_ALU_OUT_18_port, next_ALU_OUT_17_port, 
      next_ALU_OUT_16_port, next_ALU_OUT_15_port, next_ALU_OUT_14_port, 
      next_ALU_OUT_13_port, next_ALU_OUT_12_port, next_ALU_OUT_11_port, 
      next_ALU_OUT_10_port, next_ALU_OUT_9_port, next_ALU_OUT_8_port, 
      next_ALU_OUT_7_port, next_ALU_OUT_6_port, next_ALU_OUT_5_port, 
      next_ALU_OUT_4_port, next_ALU_OUT_3_port, next_ALU_OUT_2_port, 
      next_ALU_OUT_1_port, next_ALU_OUT_0_port, current_ALU_OUT_31_port, 
      current_ALU_OUT_30_port, current_ALU_OUT_29_port, current_ALU_OUT_28_port
      , current_ALU_OUT_27_port, current_ALU_OUT_26_port, 
      current_ALU_OUT_25_port, current_ALU_OUT_24_port, current_ALU_OUT_23_port
      , current_ALU_OUT_22_port, current_ALU_OUT_21_port, 
      current_ALU_OUT_20_port, current_ALU_OUT_19_port, current_ALU_OUT_18_port
      , current_ALU_OUT_17_port, current_ALU_OUT_16_port, 
      current_ALU_OUT_15_port, current_ALU_OUT_14_port, current_ALU_OUT_13_port
      , current_ALU_OUT_12_port, current_ALU_OUT_11_port, 
      current_ALU_OUT_10_port, current_ALU_OUT_9_port, current_ALU_OUT_8_port, 
      current_ALU_OUT_7_port, current_ALU_OUT_6_port, B_OUT_31_port, 
      B_OUT_30_port, B_OUT_29_port, B_OUT_28_port, B_OUT_27_port, B_OUT_26_port
      , B_OUT_25_port, B_OUT_24_port, B_OUT_23_port, B_OUT_22_port, 
      B_OUT_21_port, B_OUT_20_port, B_OUT_19_port, B_OUT_18_port, B_OUT_17_port
      , B_OUT_16_port, B_OUT_15_port, B_OUT_14_port, B_OUT_13_port, 
      B_OUT_12_port, B_OUT_11_port, B_OUT_10_port, B_OUT_9_port, B_OUT_8_port, 
      B_OUT_7_port, B_OUT_6_port, B_OUT_5_port, B_OUT_4_port, B_OUT_3_port, 
      B_OUT_2_port, B_OUT_1_port, B_OUT_0_port, current_ALU_OUT2_31_port, 
      current_ALU_OUT2_30_port, current_ALU_OUT2_29_port, 
      current_ALU_OUT2_28_port, current_ALU_OUT2_27_port, 
      current_ALU_OUT2_26_port, current_ALU_OUT2_25_port, 
      current_ALU_OUT2_24_port, current_ALU_OUT2_23_port, 
      current_ALU_OUT2_22_port, current_ALU_OUT2_21_port, 
      current_ALU_OUT2_20_port, current_ALU_OUT2_19_port, 
      current_ALU_OUT2_18_port, current_ALU_OUT2_17_port, 
      current_ALU_OUT2_16_port, current_ALU_OUT2_15_port, 
      current_ALU_OUT2_14_port, current_ALU_OUT2_13_port, 
      current_ALU_OUT2_12_port, current_ALU_OUT2_11_port, 
      current_ALU_OUT2_10_port, current_ALU_OUT2_9_port, 
      current_ALU_OUT2_8_port, current_ALU_OUT2_7_port, current_ALU_OUT2_6_port
      , current_ALU_OUT2_5_port, current_ALU_OUT2_4_port, 
      current_ALU_OUT2_3_port, current_ALU_OUT2_2_port, current_ALU_OUT2_1_port
      , current_ALU_OUT2_0_port, A_OUT_31_port, A_OUT_30_port, A_OUT_29_port, 
      A_OUT_28_port, A_OUT_27_port, A_OUT_26_port, A_OUT_25_port, A_OUT_24_port
      , A_OUT_23_port, A_OUT_22_port, A_OUT_21_port, A_OUT_20_port, 
      A_OUT_19_port, A_OUT_18_port, A_OUT_17_port, A_OUT_16_port, A_OUT_15_port
      , A_OUT_14_port, A_OUT_13_port, A_OUT_12_port, A_OUT_11_port, 
      A_OUT_10_port, A_OUT_9_port, A_OUT_8_port, A_OUT_7_port, A_OUT_6_port, 
      A_OUT_5_port, A_OUT_4_port, A_OUT_3_port, A_OUT_2_port, A_OUT_1_port, 
      A_OUT_0_port, branch_taken, PC_MUX_SEL, ALU_OP1_31_port, ALU_OP1_30_port,
      ALU_OP1_29_port, ALU_OP1_28_port, ALU_OP1_27_port, ALU_OP1_26_port, 
      ALU_OP1_25_port, ALU_OP1_24_port, ALU_OP1_23_port, ALU_OP1_22_port, 
      ALU_OP1_21_port, ALU_OP1_20_port, ALU_OP1_19_port, ALU_OP1_18_port, 
      ALU_OP1_17_port, ALU_OP1_16_port, ALU_OP1_15_port, ALU_OP1_14_port, 
      ALU_OP1_13_port, ALU_OP1_12_port, ALU_OP1_11_port, ALU_OP1_10_port, 
      ALU_OP1_9_port, ALU_OP1_8_port, ALU_OP1_7_port, ALU_OP1_6_port, 
      ALU_OP1_5_port, ALU_OP1_4_port, ALU_OP1_3_port, ALU_OP1_2_port, 
      ALU_OP1_1_port, ALU_OP1_0_port, IMM_OUT_31_port, IMM_OUT_30_port, 
      IMM_OUT_29_port, IMM_OUT_28_port, IMM_OUT_27_port, IMM_OUT_26_port, 
      IMM_OUT_25_port, IMM_OUT_24_port, IMM_OUT_23_port, IMM_OUT_22_port, 
      IMM_OUT_21_port, IMM_OUT_20_port, IMM_OUT_19_port, IMM_OUT_18_port, 
      IMM_OUT_17_port, IMM_OUT_16_port, IMM_OUT_15_port, IMM_OUT_14_port, 
      IMM_OUT_13_port, IMM_OUT_12_port, IMM_OUT_11_port, IMM_OUT_10_port, 
      IMM_OUT_9_port, IMM_OUT_8_port, IMM_OUT_7_port, IMM_OUT_6_port, 
      IMM_OUT_5_port, IMM_OUT_4_port, IMM_OUT_3_port, IMM_OUT_2_port, 
      IMM_OUT_1_port, IMM_OUT_0_port, ALU_OP2_31_port, ALU_OP2_30_port, 
      ALU_OP2_29_port, ALU_OP2_28_port, ALU_OP2_27_port, ALU_OP2_26_port, 
      ALU_OP2_25_port, ALU_OP2_24_port, ALU_OP2_23_port, ALU_OP2_22_port, 
      ALU_OP2_21_port, ALU_OP2_20_port, ALU_OP2_19_port, ALU_OP2_18_port, 
      ALU_OP2_17_port, ALU_OP2_16_port, ALU_OP2_15_port, ALU_OP2_14_port, 
      ALU_OP2_13_port, ALU_OP2_12_port, ALU_OP2_11_port, ALU_OP2_10_port, 
      ALU_OP2_9_port, ALU_OP2_8_port, ALU_OP2_7_port, ALU_OP2_6_port, 
      ALU_OP2_5_port, ALU_OP2_4_port, ALU_OP2_3_port, ALU_OP2_2_port, 
      ALU_OP2_1_port, ALU_OP2_0_port, OUT_MUX_DATA_31_port, 
      OUT_MUX_DATA_30_port, OUT_MUX_DATA_29_port, OUT_MUX_DATA_28_port, 
      OUT_MUX_DATA_27_port, OUT_MUX_DATA_26_port, OUT_MUX_DATA_25_port, 
      OUT_MUX_DATA_24_port, OUT_MUX_DATA_23_port, OUT_MUX_DATA_22_port, 
      OUT_MUX_DATA_21_port, OUT_MUX_DATA_20_port, OUT_MUX_DATA_19_port, 
      OUT_MUX_DATA_18_port, OUT_MUX_DATA_17_port, OUT_MUX_DATA_16_port, 
      OUT_MUX_DATA_15_port, OUT_MUX_DATA_14_port, OUT_MUX_DATA_13_port, 
      OUT_MUX_DATA_12_port, OUT_MUX_DATA_11_port, OUT_MUX_DATA_10_port, 
      OUT_MUX_DATA_9_port, OUT_MUX_DATA_8_port, OUT_MUX_DATA_7_port, 
      OUT_MUX_DATA_6_port, OUT_MUX_DATA_5_port, OUT_MUX_DATA_4_port, 
      OUT_MUX_DATA_3_port, OUT_MUX_DATA_2_port, OUT_MUX_DATA_1_port, 
      OUT_MUX_DATA_0_port, WB_DATA_31_port, WB_DATA_30_port, WB_DATA_29_port, 
      WB_DATA_28_port, WB_DATA_27_port, WB_DATA_26_port, WB_DATA_25_port, 
      WB_DATA_24_port, WB_DATA_23_port, WB_DATA_22_port, WB_DATA_21_port, 
      WB_DATA_20_port, WB_DATA_19_port, WB_DATA_18_port, WB_DATA_17_port, 
      WB_DATA_16_port, WB_DATA_15_port, WB_DATA_14_port, WB_DATA_13_port, 
      WB_DATA_12_port, WB_DATA_11_port, WB_DATA_10_port, WB_DATA_9_port, 
      WB_DATA_8_port, WB_DATA_7_port, WB_DATA_6_port, WB_DATA_5_port, 
      WB_DATA_4_port, WB_DATA_3_port, WB_DATA_2_port, WB_DATA_1_port, 
      WB_DATA_0_port, WB_ADDR_4_port, WB_ADDR_3_port, WB_ADDR_2_port, 
      WB_ADDR_1_port, WB_ADDR_0_port, n_2152, n_2153, n_2154, n_2155, n_2156, 
      n_2157 : std_logic;

begin
   D_ADDR <= ( D_ADDR_5_port, D_ADDR_4_port, D_ADDR_3_port, D_ADDR_2_port, 
      D_ADDR_1_port, D_ADDR_0_port );
   PC_BUS <= ( PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port );
   
   RF : REGISTER_FILE_NBIT32_NREG32 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, RD1 => RegA_LATCH_EN, RD2 => 
                           RegB_LATCH_EN, WR => RF_WE, ADD_WR(4) => 
                           WB_ADDR_4_port, ADD_WR(3) => WB_ADDR_3_port, 
                           ADD_WR(2) => WB_ADDR_2_port, ADD_WR(1) => 
                           WB_ADDR_1_port, ADD_WR(0) => WB_ADDR_0_port, 
                           ADD_RD1(4) => current_IW_25_port, ADD_RD1(3) => 
                           current_IW_24_port, ADD_RD1(2) => current_IW_23_port
                           , ADD_RD1(1) => current_IW_22_port, ADD_RD1(0) => 
                           current_IW_21_port, ADD_RD2(4) => current_IW_20_port
                           , ADD_RD2(3) => current_IW_19_port, ADD_RD2(2) => 
                           current_IW_18_port, ADD_RD2(1) => current_IW_17_port
                           , ADD_RD2(0) => current_IW_16_port, DATAIN(31) => 
                           WB_DATA_31_port, DATAIN(30) => WB_DATA_30_port, 
                           DATAIN(29) => WB_DATA_29_port, DATAIN(28) => 
                           WB_DATA_28_port, DATAIN(27) => WB_DATA_27_port, 
                           DATAIN(26) => WB_DATA_26_port, DATAIN(25) => 
                           WB_DATA_25_port, DATAIN(24) => WB_DATA_24_port, 
                           DATAIN(23) => WB_DATA_23_port, DATAIN(22) => 
                           WB_DATA_22_port, DATAIN(21) => WB_DATA_21_port, 
                           DATAIN(20) => WB_DATA_20_port, DATAIN(19) => 
                           WB_DATA_19_port, DATAIN(18) => WB_DATA_18_port, 
                           DATAIN(17) => WB_DATA_17_port, DATAIN(16) => 
                           WB_DATA_16_port, DATAIN(15) => WB_DATA_15_port, 
                           DATAIN(14) => WB_DATA_14_port, DATAIN(13) => 
                           WB_DATA_13_port, DATAIN(12) => WB_DATA_12_port, 
                           DATAIN(11) => WB_DATA_11_port, DATAIN(10) => 
                           WB_DATA_10_port, DATAIN(9) => WB_DATA_9_port, 
                           DATAIN(8) => WB_DATA_8_port, DATAIN(7) => 
                           WB_DATA_7_port, DATAIN(6) => WB_DATA_6_port, 
                           DATAIN(5) => WB_DATA_5_port, DATAIN(4) => 
                           WB_DATA_4_port, DATAIN(3) => WB_DATA_3_port, 
                           DATAIN(2) => WB_DATA_2_port, DATAIN(1) => 
                           WB_DATA_1_port, DATAIN(0) => WB_DATA_0_port, 
                           OUT1(31) => A_OUT_31_port, OUT1(30) => A_OUT_30_port
                           , OUT1(29) => A_OUT_29_port, OUT1(28) => 
                           A_OUT_28_port, OUT1(27) => A_OUT_27_port, OUT1(26) 
                           => A_OUT_26_port, OUT1(25) => A_OUT_25_port, 
                           OUT1(24) => A_OUT_24_port, OUT1(23) => A_OUT_23_port
                           , OUT1(22) => A_OUT_22_port, OUT1(21) => 
                           A_OUT_21_port, OUT1(20) => A_OUT_20_port, OUT1(19) 
                           => A_OUT_19_port, OUT1(18) => A_OUT_18_port, 
                           OUT1(17) => A_OUT_17_port, OUT1(16) => A_OUT_16_port
                           , OUT1(15) => A_OUT_15_port, OUT1(14) => 
                           A_OUT_14_port, OUT1(13) => A_OUT_13_port, OUT1(12) 
                           => A_OUT_12_port, OUT1(11) => A_OUT_11_port, 
                           OUT1(10) => A_OUT_10_port, OUT1(9) => A_OUT_9_port, 
                           OUT1(8) => A_OUT_8_port, OUT1(7) => A_OUT_7_port, 
                           OUT1(6) => A_OUT_6_port, OUT1(5) => A_OUT_5_port, 
                           OUT1(4) => A_OUT_4_port, OUT1(3) => A_OUT_3_port, 
                           OUT1(2) => A_OUT_2_port, OUT1(1) => A_OUT_1_port, 
                           OUT1(0) => A_OUT_0_port, OUT2(31) => B_OUT_31_port, 
                           OUT2(30) => B_OUT_30_port, OUT2(29) => B_OUT_29_port
                           , OUT2(28) => B_OUT_28_port, OUT2(27) => 
                           B_OUT_27_port, OUT2(26) => B_OUT_26_port, OUT2(25) 
                           => B_OUT_25_port, OUT2(24) => B_OUT_24_port, 
                           OUT2(23) => B_OUT_23_port, OUT2(22) => B_OUT_22_port
                           , OUT2(21) => B_OUT_21_port, OUT2(20) => 
                           B_OUT_20_port, OUT2(19) => B_OUT_19_port, OUT2(18) 
                           => B_OUT_18_port, OUT2(17) => B_OUT_17_port, 
                           OUT2(16) => B_OUT_16_port, OUT2(15) => B_OUT_15_port
                           , OUT2(14) => B_OUT_14_port, OUT2(13) => 
                           B_OUT_13_port, OUT2(12) => B_OUT_12_port, OUT2(11) 
                           => B_OUT_11_port, OUT2(10) => B_OUT_10_port, OUT2(9)
                           => B_OUT_9_port, OUT2(8) => B_OUT_8_port, OUT2(7) =>
                           B_OUT_7_port, OUT2(6) => B_OUT_6_port, OUT2(5) => 
                           B_OUT_5_port, OUT2(4) => B_OUT_4_port, OUT2(3) => 
                           B_OUT_3_port, OUT2(2) => B_OUT_2_port, OUT2(1) => 
                           B_OUT_1_port, OUT2(0) => B_OUT_0_port);
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   PC_REG : REG_GENERIC_NBIT32_8 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => PC_IN(31), DATA_IN(30) 
                           => PC_IN(30), DATA_IN(29) => PC_IN(29), DATA_IN(28) 
                           => PC_IN(28), DATA_IN(27) => PC_IN(27), DATA_IN(26) 
                           => PC_IN(26), DATA_IN(25) => PC_IN(25), DATA_IN(24) 
                           => PC_IN(24), DATA_IN(23) => PC_IN(23), DATA_IN(22) 
                           => PC_IN(22), DATA_IN(21) => PC_IN(21), DATA_IN(20) 
                           => PC_IN(20), DATA_IN(19) => PC_IN(19), DATA_IN(18) 
                           => PC_IN(18), DATA_IN(17) => PC_IN(17), DATA_IN(16) 
                           => PC_IN(16), DATA_IN(15) => PC_IN(15), DATA_IN(14) 
                           => PC_IN(14), DATA_IN(13) => PC_IN(13), DATA_IN(12) 
                           => PC_IN(12), DATA_IN(11) => PC_IN(11), DATA_IN(10) 
                           => PC_IN(10), DATA_IN(9) => PC_IN(9), DATA_IN(8) => 
                           PC_IN(8), DATA_IN(7) => PC_IN(7), DATA_IN(6) => 
                           PC_IN(6), DATA_IN(5) => PC_IN(5), DATA_IN(4) => 
                           PC_IN(4), DATA_IN(3) => PC_IN(3), DATA_IN(2) => 
                           PC_IN(2), DATA_IN(1) => PC_IN(1), DATA_IN(0) => 
                           PC_IN(0), DATA_OUT(31) => current_PC1_31_port, 
                           DATA_OUT(30) => current_PC1_30_port, DATA_OUT(29) =>
                           current_PC1_29_port, DATA_OUT(28) => 
                           current_PC1_28_port, DATA_OUT(27) => 
                           current_PC1_27_port, DATA_OUT(26) => 
                           current_PC1_26_port, DATA_OUT(25) => 
                           current_PC1_25_port, DATA_OUT(24) => 
                           current_PC1_24_port, DATA_OUT(23) => 
                           current_PC1_23_port, DATA_OUT(22) => 
                           current_PC1_22_port, DATA_OUT(21) => 
                           current_PC1_21_port, DATA_OUT(20) => 
                           current_PC1_20_port, DATA_OUT(19) => 
                           current_PC1_19_port, DATA_OUT(18) => 
                           current_PC1_18_port, DATA_OUT(17) => 
                           current_PC1_17_port, DATA_OUT(16) => 
                           current_PC1_16_port, DATA_OUT(15) => 
                           current_PC1_15_port, DATA_OUT(14) => 
                           current_PC1_14_port, DATA_OUT(13) => 
                           current_PC1_13_port, DATA_OUT(12) => 
                           current_PC1_12_port, DATA_OUT(11) => 
                           current_PC1_11_port, DATA_OUT(10) => 
                           current_PC1_10_port, DATA_OUT(9) => 
                           current_PC1_9_port, DATA_OUT(8) => 
                           current_PC1_8_port, DATA_OUT(7) => 
                           current_PC1_7_port, DATA_OUT(6) => 
                           current_PC1_6_port, DATA_OUT(5) => 
                           current_PC1_5_port, DATA_OUT(4) => 
                           current_PC1_4_port, DATA_OUT(3) => 
                           current_PC1_3_port, DATA_OUT(2) => 
                           current_PC1_2_port, DATA_OUT(1) => 
                           current_PC1_1_port, DATA_OUT(0) => 
                           current_PC1_0_port);
   PC2_REG : REG_GENERIC_NBIT32_7 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => current_PC1_31_port, 
                           DATA_IN(30) => current_PC1_30_port, DATA_IN(29) => 
                           current_PC1_29_port, DATA_IN(28) => 
                           current_PC1_28_port, DATA_IN(27) => 
                           current_PC1_27_port, DATA_IN(26) => 
                           current_PC1_26_port, DATA_IN(25) => 
                           current_PC1_25_port, DATA_IN(24) => 
                           current_PC1_24_port, DATA_IN(23) => 
                           current_PC1_23_port, DATA_IN(22) => 
                           current_PC1_22_port, DATA_IN(21) => 
                           current_PC1_21_port, DATA_IN(20) => 
                           current_PC1_20_port, DATA_IN(19) => 
                           current_PC1_19_port, DATA_IN(18) => 
                           current_PC1_18_port, DATA_IN(17) => 
                           current_PC1_17_port, DATA_IN(16) => 
                           current_PC1_16_port, DATA_IN(15) => 
                           current_PC1_15_port, DATA_IN(14) => 
                           current_PC1_14_port, DATA_IN(13) => 
                           current_PC1_13_port, DATA_IN(12) => 
                           current_PC1_12_port, DATA_IN(11) => 
                           current_PC1_11_port, DATA_IN(10) => 
                           current_PC1_10_port, DATA_IN(9) => 
                           current_PC1_9_port, DATA_IN(8) => current_PC1_8_port
                           , DATA_IN(7) => current_PC1_7_port, DATA_IN(6) => 
                           current_PC1_6_port, DATA_IN(5) => current_PC1_5_port
                           , DATA_IN(4) => current_PC1_4_port, DATA_IN(3) => 
                           current_PC1_3_port, DATA_IN(2) => current_PC1_2_port
                           , DATA_IN(1) => current_PC1_1_port, DATA_IN(0) => 
                           current_PC1_0_port, DATA_OUT(31) => 
                           current_PC2_31_port, DATA_OUT(30) => 
                           current_PC2_30_port, DATA_OUT(29) => 
                           current_PC2_29_port, DATA_OUT(28) => 
                           current_PC2_28_port, DATA_OUT(27) => 
                           current_PC2_27_port, DATA_OUT(26) => 
                           current_PC2_26_port, DATA_OUT(25) => 
                           current_PC2_25_port, DATA_OUT(24) => 
                           current_PC2_24_port, DATA_OUT(23) => 
                           current_PC2_23_port, DATA_OUT(22) => 
                           current_PC2_22_port, DATA_OUT(21) => 
                           current_PC2_21_port, DATA_OUT(20) => 
                           current_PC2_20_port, DATA_OUT(19) => 
                           current_PC2_19_port, DATA_OUT(18) => 
                           current_PC2_18_port, DATA_OUT(17) => 
                           current_PC2_17_port, DATA_OUT(16) => 
                           current_PC2_16_port, DATA_OUT(15) => 
                           current_PC2_15_port, DATA_OUT(14) => 
                           current_PC2_14_port, DATA_OUT(13) => 
                           current_PC2_13_port, DATA_OUT(12) => 
                           current_PC2_12_port, DATA_OUT(11) => 
                           current_PC2_11_port, DATA_OUT(10) => 
                           current_PC2_10_port, DATA_OUT(9) => 
                           current_PC2_9_port, DATA_OUT(8) => 
                           current_PC2_8_port, DATA_OUT(7) => 
                           current_PC2_7_port, DATA_OUT(6) => 
                           current_PC2_6_port, DATA_OUT(5) => 
                           current_PC2_5_port, DATA_OUT(4) => 
                           current_PC2_4_port, DATA_OUT(3) => 
                           current_PC2_3_port, DATA_OUT(2) => 
                           current_PC2_2_port, DATA_OUT(1) => 
                           current_PC2_1_port, DATA_OUT(0) => 
                           current_PC2_0_port);
   PC3_REG : REG_GENERIC_NBIT32_6 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => current_PC2_31_port, 
                           DATA_IN(30) => current_PC2_30_port, DATA_IN(29) => 
                           current_PC2_29_port, DATA_IN(28) => 
                           current_PC2_28_port, DATA_IN(27) => 
                           current_PC2_27_port, DATA_IN(26) => 
                           current_PC2_26_port, DATA_IN(25) => 
                           current_PC2_25_port, DATA_IN(24) => 
                           current_PC2_24_port, DATA_IN(23) => 
                           current_PC2_23_port, DATA_IN(22) => 
                           current_PC2_22_port, DATA_IN(21) => 
                           current_PC2_21_port, DATA_IN(20) => 
                           current_PC2_20_port, DATA_IN(19) => 
                           current_PC2_19_port, DATA_IN(18) => 
                           current_PC2_18_port, DATA_IN(17) => 
                           current_PC2_17_port, DATA_IN(16) => 
                           current_PC2_16_port, DATA_IN(15) => 
                           current_PC2_15_port, DATA_IN(14) => 
                           current_PC2_14_port, DATA_IN(13) => 
                           current_PC2_13_port, DATA_IN(12) => 
                           current_PC2_12_port, DATA_IN(11) => 
                           current_PC2_11_port, DATA_IN(10) => 
                           current_PC2_10_port, DATA_IN(9) => 
                           current_PC2_9_port, DATA_IN(8) => current_PC2_8_port
                           , DATA_IN(7) => current_PC2_7_port, DATA_IN(6) => 
                           current_PC2_6_port, DATA_IN(5) => current_PC2_5_port
                           , DATA_IN(4) => current_PC2_4_port, DATA_IN(3) => 
                           current_PC2_3_port, DATA_IN(2) => current_PC2_2_port
                           , DATA_IN(1) => current_PC2_1_port, DATA_IN(0) => 
                           current_PC2_0_port, DATA_OUT(31) => 
                           current_PC3_31_port, DATA_OUT(30) => 
                           current_PC3_30_port, DATA_OUT(29) => 
                           current_PC3_29_port, DATA_OUT(28) => 
                           current_PC3_28_port, DATA_OUT(27) => 
                           current_PC3_27_port, DATA_OUT(26) => 
                           current_PC3_26_port, DATA_OUT(25) => 
                           current_PC3_25_port, DATA_OUT(24) => 
                           current_PC3_24_port, DATA_OUT(23) => 
                           current_PC3_23_port, DATA_OUT(22) => 
                           current_PC3_22_port, DATA_OUT(21) => 
                           current_PC3_21_port, DATA_OUT(20) => 
                           current_PC3_20_port, DATA_OUT(19) => 
                           current_PC3_19_port, DATA_OUT(18) => 
                           current_PC3_18_port, DATA_OUT(17) => 
                           current_PC3_17_port, DATA_OUT(16) => 
                           current_PC3_16_port, DATA_OUT(15) => 
                           current_PC3_15_port, DATA_OUT(14) => 
                           current_PC3_14_port, DATA_OUT(13) => 
                           current_PC3_13_port, DATA_OUT(12) => 
                           current_PC3_12_port, DATA_OUT(11) => 
                           current_PC3_11_port, DATA_OUT(10) => 
                           current_PC3_10_port, DATA_OUT(9) => 
                           current_PC3_9_port, DATA_OUT(8) => 
                           current_PC3_8_port, DATA_OUT(7) => 
                           current_PC3_7_port, DATA_OUT(6) => 
                           current_PC3_6_port, DATA_OUT(5) => 
                           current_PC3_5_port, DATA_OUT(4) => 
                           current_PC3_4_port, DATA_OUT(3) => 
                           current_PC3_3_port, DATA_OUT(2) => 
                           current_PC3_2_port, DATA_OUT(1) => 
                           current_PC3_1_port, DATA_OUT(0) => 
                           current_PC3_0_port);
   NPC_REG : REG_GENERIC_NBIT32_5 port map( CLK => CLK, RST => RST, EN => 
                           NPC_LATCH_EN, DATA_IN(31) => next_NPC_31_port, 
                           DATA_IN(30) => next_NPC_30_port, DATA_IN(29) => 
                           next_NPC_29_port, DATA_IN(28) => next_NPC_28_port, 
                           DATA_IN(27) => next_NPC_27_port, DATA_IN(26) => 
                           next_NPC_26_port, DATA_IN(25) => next_NPC_25_port, 
                           DATA_IN(24) => next_NPC_24_port, DATA_IN(23) => 
                           next_NPC_23_port, DATA_IN(22) => next_NPC_22_port, 
                           DATA_IN(21) => next_NPC_21_port, DATA_IN(20) => 
                           next_NPC_20_port, DATA_IN(19) => next_NPC_19_port, 
                           DATA_IN(18) => next_NPC_18_port, DATA_IN(17) => 
                           next_NPC_17_port, DATA_IN(16) => next_NPC_16_port, 
                           DATA_IN(15) => next_NPC_15_port, DATA_IN(14) => 
                           next_NPC_14_port, DATA_IN(13) => next_NPC_13_port, 
                           DATA_IN(12) => next_NPC_12_port, DATA_IN(11) => 
                           next_NPC_11_port, DATA_IN(10) => next_NPC_10_port, 
                           DATA_IN(9) => next_NPC_9_port, DATA_IN(8) => 
                           next_NPC_8_port, DATA_IN(7) => next_NPC_7_port, 
                           DATA_IN(6) => next_NPC_6_port, DATA_IN(5) => 
                           next_NPC_5_port, DATA_IN(4) => next_NPC_4_port, 
                           DATA_IN(3) => next_NPC_3_port, DATA_IN(2) => 
                           next_NPC_2_port, DATA_IN(1) => next_NPC_1_port, 
                           DATA_IN(0) => next_NPC_0_port, DATA_OUT(31) => 
                           current_NPC_31_port, DATA_OUT(30) => 
                           current_NPC_30_port, DATA_OUT(29) => 
                           current_NPC_29_port, DATA_OUT(28) => 
                           current_NPC_28_port, DATA_OUT(27) => 
                           current_NPC_27_port, DATA_OUT(26) => 
                           current_NPC_26_port, DATA_OUT(25) => 
                           current_NPC_25_port, DATA_OUT(24) => 
                           current_NPC_24_port, DATA_OUT(23) => 
                           current_NPC_23_port, DATA_OUT(22) => 
                           current_NPC_22_port, DATA_OUT(21) => 
                           current_NPC_21_port, DATA_OUT(20) => 
                           current_NPC_20_port, DATA_OUT(19) => 
                           current_NPC_19_port, DATA_OUT(18) => 
                           current_NPC_18_port, DATA_OUT(17) => 
                           current_NPC_17_port, DATA_OUT(16) => 
                           current_NPC_16_port, DATA_OUT(15) => 
                           current_NPC_15_port, DATA_OUT(14) => 
                           current_NPC_14_port, DATA_OUT(13) => 
                           current_NPC_13_port, DATA_OUT(12) => 
                           current_NPC_12_port, DATA_OUT(11) => 
                           current_NPC_11_port, DATA_OUT(10) => 
                           current_NPC_10_port, DATA_OUT(9) => 
                           current_NPC_9_port, DATA_OUT(8) => 
                           current_NPC_8_port, DATA_OUT(7) => 
                           current_NPC_7_port, DATA_OUT(6) => 
                           current_NPC_6_port, DATA_OUT(5) => 
                           current_NPC_5_port, DATA_OUT(4) => 
                           current_NPC_4_port, DATA_OUT(3) => 
                           current_NPC_3_port, DATA_OUT(2) => 
                           current_NPC_2_port, DATA_OUT(1) => 
                           current_NPC_1_port, DATA_OUT(0) => 
                           current_NPC_0_port);
   IR_REG : REG_GENERIC_NBIT32_4 port map( CLK => CLK, RST => RST, EN => 
                           IR_LATCH_EN, DATA_IN(31) => IR_IN(31), DATA_IN(30) 
                           => IR_IN(30), DATA_IN(29) => IR_IN(29), DATA_IN(28) 
                           => IR_IN(28), DATA_IN(27) => IR_IN(27), DATA_IN(26) 
                           => IR_IN(26), DATA_IN(25) => IR_IN(25), DATA_IN(24) 
                           => IR_IN(24), DATA_IN(23) => IR_IN(23), DATA_IN(22) 
                           => IR_IN(22), DATA_IN(21) => IR_IN(21), DATA_IN(20) 
                           => IR_IN(20), DATA_IN(19) => IR_IN(19), DATA_IN(18) 
                           => IR_IN(18), DATA_IN(17) => IR_IN(17), DATA_IN(16) 
                           => IR_IN(16), DATA_IN(15) => IR_IN(15), DATA_IN(14) 
                           => IR_IN(14), DATA_IN(13) => IR_IN(13), DATA_IN(12) 
                           => IR_IN(12), DATA_IN(11) => IR_IN(11), DATA_IN(10) 
                           => IR_IN(10), DATA_IN(9) => IR_IN(9), DATA_IN(8) => 
                           IR_IN(8), DATA_IN(7) => IR_IN(7), DATA_IN(6) => 
                           IR_IN(6), DATA_IN(5) => IR_IN(5), DATA_IN(4) => 
                           IR_IN(4), DATA_IN(3) => IR_IN(3), DATA_IN(2) => 
                           IR_IN(2), DATA_IN(1) => IR_IN(1), DATA_IN(0) => 
                           IR_IN(0), DATA_OUT(31) => n_2152, DATA_OUT(30) => 
                           n_2153, DATA_OUT(29) => n_2154, DATA_OUT(28) => 
                           n_2155, DATA_OUT(27) => n_2156, DATA_OUT(26) => 
                           n_2157, DATA_OUT(25) => current_IW_25_port, 
                           DATA_OUT(24) => current_IW_24_port, DATA_OUT(23) => 
                           current_IW_23_port, DATA_OUT(22) => 
                           current_IW_22_port, DATA_OUT(21) => 
                           current_IW_21_port, DATA_OUT(20) => 
                           current_IW_20_port, DATA_OUT(19) => 
                           current_IW_19_port, DATA_OUT(18) => 
                           current_IW_18_port, DATA_OUT(17) => 
                           current_IW_17_port, DATA_OUT(16) => 
                           current_IW_16_port, DATA_OUT(15) => 
                           current_IW_15_port, DATA_OUT(14) => 
                           current_IW_14_port, DATA_OUT(13) => 
                           current_IW_13_port, DATA_OUT(12) => 
                           current_IW_12_port, DATA_OUT(11) => 
                           current_IW_11_port, DATA_OUT(10) => 
                           current_IW_10_port, DATA_OUT(9) => current_IW_9_port
                           , DATA_OUT(8) => current_IW_8_port, DATA_OUT(7) => 
                           current_IW_7_port, DATA_OUT(6) => current_IW_6_port,
                           DATA_OUT(5) => current_IW_5_port, DATA_OUT(4) => 
                           current_IW_4_port, DATA_OUT(3) => current_IW_3_port,
                           DATA_OUT(2) => current_IW_2_port, DATA_OUT(1) => 
                           current_IW_1_port, DATA_OUT(0) => current_IW_0_port)
                           ;
   IMM_REG : REG_GENERIC_NBIT16 port map( CLK => CLK, RST => RST, EN => 
                           RegIMM_LATCH_EN, DATA_IN(15) => current_IW_15_port, 
                           DATA_IN(14) => current_IW_14_port, DATA_IN(13) => 
                           current_IW_13_port, DATA_IN(12) => 
                           current_IW_12_port, DATA_IN(11) => 
                           current_IW_11_port, DATA_IN(10) => 
                           current_IW_10_port, DATA_IN(9) => current_IW_9_port,
                           DATA_IN(8) => current_IW_8_port, DATA_IN(7) => 
                           current_IW_7_port, DATA_IN(6) => current_IW_6_port, 
                           DATA_IN(5) => current_IW_5_port, DATA_IN(4) => 
                           current_IW_4_port, DATA_IN(3) => current_IW_3_port, 
                           DATA_IN(2) => current_IW_2_port, DATA_IN(1) => 
                           current_IW_1_port, DATA_IN(0) => current_IW_0_port, 
                           DATA_OUT(15) => IMM_IN_15_port, DATA_OUT(14) => 
                           IMM_IN_14_port, DATA_OUT(13) => IMM_IN_13_port, 
                           DATA_OUT(12) => IMM_IN_12_port, DATA_OUT(11) => 
                           IMM_IN_11_port, DATA_OUT(10) => IMM_IN_10_port, 
                           DATA_OUT(9) => IMM_IN_9_port, DATA_OUT(8) => 
                           IMM_IN_8_port, DATA_OUT(7) => IMM_IN_7_port, 
                           DATA_OUT(6) => IMM_IN_6_port, DATA_OUT(5) => 
                           IMM_IN_5_port, DATA_OUT(4) => IMM_IN_4_port, 
                           DATA_OUT(3) => IMM_IN_3_port, DATA_OUT(2) => 
                           IMM_IN_2_port, DATA_OUT(1) => IMM_IN_1_port, 
                           DATA_OUT(0) => IMM_IN_0_port);
   WB1_REG : REG_GENERIC_NBIT5_0 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, DATA_IN(4) => WB1_IN_4_port, 
                           DATA_IN(3) => WB1_IN_3_port, DATA_IN(2) => 
                           WB1_IN_2_port, DATA_IN(1) => WB1_IN_1_port, 
                           DATA_IN(0) => WB1_IN_0_port, DATA_OUT(4) => 
                           WB2_IN_4_port, DATA_OUT(3) => WB2_IN_3_port, 
                           DATA_OUT(2) => WB2_IN_2_port, DATA_OUT(1) => 
                           WB2_IN_1_port, DATA_OUT(0) => WB2_IN_0_port);
   WB2_REG : REG_GENERIC_NBIT5_2 port map( CLK => CLK, RST => RST, EN => 
                           ALU_OUTREG_EN, DATA_IN(4) => WB2_IN_4_port, 
                           DATA_IN(3) => WB2_IN_3_port, DATA_IN(2) => 
                           WB2_IN_2_port, DATA_IN(1) => WB2_IN_1_port, 
                           DATA_IN(0) => WB2_IN_0_port, DATA_OUT(4) => 
                           WB2_OUT_4_port, DATA_OUT(3) => WB2_OUT_3_port, 
                           DATA_OUT(2) => WB2_OUT_2_port, DATA_OUT(1) => 
                           WB2_OUT_1_port, DATA_OUT(0) => WB2_OUT_0_port);
   WB3_REG : REG_GENERIC_NBIT5_1 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, DATA_IN(4) => WB2_OUT_4_port, 
                           DATA_IN(3) => WB2_OUT_3_port, DATA_IN(2) => 
                           WB2_OUT_2_port, DATA_IN(1) => WB2_OUT_1_port, 
                           DATA_IN(0) => WB2_OUT_0_port, DATA_OUT(4) => 
                           WB3_OUT_4_port, DATA_OUT(3) => WB3_OUT_3_port, 
                           DATA_OUT(2) => WB3_OUT_2_port, DATA_OUT(1) => 
                           WB3_OUT_1_port, DATA_OUT(0) => WB3_OUT_0_port);
   ALU_OUT_REG : REG_GENERIC_NBIT32_3 port map( CLK => CLK, RST => RST, EN => 
                           ALU_OUTREG_EN, DATA_IN(31) => next_ALU_OUT_31_port, 
                           DATA_IN(30) => next_ALU_OUT_30_port, DATA_IN(29) => 
                           next_ALU_OUT_29_port, DATA_IN(28) => 
                           next_ALU_OUT_28_port, DATA_IN(27) => 
                           next_ALU_OUT_27_port, DATA_IN(26) => 
                           next_ALU_OUT_26_port, DATA_IN(25) => 
                           next_ALU_OUT_25_port, DATA_IN(24) => 
                           next_ALU_OUT_24_port, DATA_IN(23) => 
                           next_ALU_OUT_23_port, DATA_IN(22) => 
                           next_ALU_OUT_22_port, DATA_IN(21) => 
                           next_ALU_OUT_21_port, DATA_IN(20) => 
                           next_ALU_OUT_20_port, DATA_IN(19) => 
                           next_ALU_OUT_19_port, DATA_IN(18) => 
                           next_ALU_OUT_18_port, DATA_IN(17) => 
                           next_ALU_OUT_17_port, DATA_IN(16) => 
                           next_ALU_OUT_16_port, DATA_IN(15) => 
                           next_ALU_OUT_15_port, DATA_IN(14) => 
                           next_ALU_OUT_14_port, DATA_IN(13) => 
                           next_ALU_OUT_13_port, DATA_IN(12) => 
                           next_ALU_OUT_12_port, DATA_IN(11) => 
                           next_ALU_OUT_11_port, DATA_IN(10) => 
                           next_ALU_OUT_10_port, DATA_IN(9) => 
                           next_ALU_OUT_9_port, DATA_IN(8) => 
                           next_ALU_OUT_8_port, DATA_IN(7) => 
                           next_ALU_OUT_7_port, DATA_IN(6) => 
                           next_ALU_OUT_6_port, DATA_IN(5) => 
                           next_ALU_OUT_5_port, DATA_IN(4) => 
                           next_ALU_OUT_4_port, DATA_IN(3) => 
                           next_ALU_OUT_3_port, DATA_IN(2) => 
                           next_ALU_OUT_2_port, DATA_IN(1) => 
                           next_ALU_OUT_1_port, DATA_IN(0) => 
                           next_ALU_OUT_0_port, DATA_OUT(31) => 
                           current_ALU_OUT_31_port, DATA_OUT(30) => 
                           current_ALU_OUT_30_port, DATA_OUT(29) => 
                           current_ALU_OUT_29_port, DATA_OUT(28) => 
                           current_ALU_OUT_28_port, DATA_OUT(27) => 
                           current_ALU_OUT_27_port, DATA_OUT(26) => 
                           current_ALU_OUT_26_port, DATA_OUT(25) => 
                           current_ALU_OUT_25_port, DATA_OUT(24) => 
                           current_ALU_OUT_24_port, DATA_OUT(23) => 
                           current_ALU_OUT_23_port, DATA_OUT(22) => 
                           current_ALU_OUT_22_port, DATA_OUT(21) => 
                           current_ALU_OUT_21_port, DATA_OUT(20) => 
                           current_ALU_OUT_20_port, DATA_OUT(19) => 
                           current_ALU_OUT_19_port, DATA_OUT(18) => 
                           current_ALU_OUT_18_port, DATA_OUT(17) => 
                           current_ALU_OUT_17_port, DATA_OUT(16) => 
                           current_ALU_OUT_16_port, DATA_OUT(15) => 
                           current_ALU_OUT_15_port, DATA_OUT(14) => 
                           current_ALU_OUT_14_port, DATA_OUT(13) => 
                           current_ALU_OUT_13_port, DATA_OUT(12) => 
                           current_ALU_OUT_12_port, DATA_OUT(11) => 
                           current_ALU_OUT_11_port, DATA_OUT(10) => 
                           current_ALU_OUT_10_port, DATA_OUT(9) => 
                           current_ALU_OUT_9_port, DATA_OUT(8) => 
                           current_ALU_OUT_8_port, DATA_OUT(7) => 
                           current_ALU_OUT_7_port, DATA_OUT(6) => 
                           current_ALU_OUT_6_port, DATA_OUT(5) => D_ADDR_5_port
                           , DATA_OUT(4) => D_ADDR_4_port, DATA_OUT(3) => 
                           D_ADDR_3_port, DATA_OUT(2) => D_ADDR_2_port, 
                           DATA_OUT(1) => D_ADDR_1_port, DATA_OUT(0) => 
                           D_ADDR_0_port);
   B_OUT_REG : REG_GENERIC_NBIT32_2 port map( CLK => CLK, RST => RST, EN => 
                           ALU_OUTREG_EN, DATA_IN(31) => B_OUT_31_port, 
                           DATA_IN(30) => B_OUT_30_port, DATA_IN(29) => 
                           B_OUT_29_port, DATA_IN(28) => B_OUT_28_port, 
                           DATA_IN(27) => B_OUT_27_port, DATA_IN(26) => 
                           B_OUT_26_port, DATA_IN(25) => B_OUT_25_port, 
                           DATA_IN(24) => B_OUT_24_port, DATA_IN(23) => 
                           B_OUT_23_port, DATA_IN(22) => B_OUT_22_port, 
                           DATA_IN(21) => B_OUT_21_port, DATA_IN(20) => 
                           B_OUT_20_port, DATA_IN(19) => B_OUT_19_port, 
                           DATA_IN(18) => B_OUT_18_port, DATA_IN(17) => 
                           B_OUT_17_port, DATA_IN(16) => B_OUT_16_port, 
                           DATA_IN(15) => B_OUT_15_port, DATA_IN(14) => 
                           B_OUT_14_port, DATA_IN(13) => B_OUT_13_port, 
                           DATA_IN(12) => B_OUT_12_port, DATA_IN(11) => 
                           B_OUT_11_port, DATA_IN(10) => B_OUT_10_port, 
                           DATA_IN(9) => B_OUT_9_port, DATA_IN(8) => 
                           B_OUT_8_port, DATA_IN(7) => B_OUT_7_port, DATA_IN(6)
                           => B_OUT_6_port, DATA_IN(5) => B_OUT_5_port, 
                           DATA_IN(4) => B_OUT_4_port, DATA_IN(3) => 
                           B_OUT_3_port, DATA_IN(2) => B_OUT_2_port, DATA_IN(1)
                           => B_OUT_1_port, DATA_IN(0) => B_OUT_0_port, 
                           DATA_OUT(31) => D_DATA_IN(31), DATA_OUT(30) => 
                           D_DATA_IN(30), DATA_OUT(29) => D_DATA_IN(29), 
                           DATA_OUT(28) => D_DATA_IN(28), DATA_OUT(27) => 
                           D_DATA_IN(27), DATA_OUT(26) => D_DATA_IN(26), 
                           DATA_OUT(25) => D_DATA_IN(25), DATA_OUT(24) => 
                           D_DATA_IN(24), DATA_OUT(23) => D_DATA_IN(23), 
                           DATA_OUT(22) => D_DATA_IN(22), DATA_OUT(21) => 
                           D_DATA_IN(21), DATA_OUT(20) => D_DATA_IN(20), 
                           DATA_OUT(19) => D_DATA_IN(19), DATA_OUT(18) => 
                           D_DATA_IN(18), DATA_OUT(17) => D_DATA_IN(17), 
                           DATA_OUT(16) => D_DATA_IN(16), DATA_OUT(15) => 
                           D_DATA_IN(15), DATA_OUT(14) => D_DATA_IN(14), 
                           DATA_OUT(13) => D_DATA_IN(13), DATA_OUT(12) => 
                           D_DATA_IN(12), DATA_OUT(11) => D_DATA_IN(11), 
                           DATA_OUT(10) => D_DATA_IN(10), DATA_OUT(9) => 
                           D_DATA_IN(9), DATA_OUT(8) => D_DATA_IN(8), 
                           DATA_OUT(7) => D_DATA_IN(7), DATA_OUT(6) => 
                           D_DATA_IN(6), DATA_OUT(5) => D_DATA_IN(5), 
                           DATA_OUT(4) => D_DATA_IN(4), DATA_OUT(3) => 
                           D_DATA_IN(3), DATA_OUT(2) => D_DATA_IN(2), 
                           DATA_OUT(1) => D_DATA_IN(1), DATA_OUT(0) => 
                           D_DATA_IN(0));
   ALU_OUT_REG2 : REG_GENERIC_NBIT32_1 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, DATA_IN(31) => 
                           current_ALU_OUT_31_port, DATA_IN(30) => 
                           current_ALU_OUT_30_port, DATA_IN(29) => 
                           current_ALU_OUT_29_port, DATA_IN(28) => 
                           current_ALU_OUT_28_port, DATA_IN(27) => 
                           current_ALU_OUT_27_port, DATA_IN(26) => 
                           current_ALU_OUT_26_port, DATA_IN(25) => 
                           current_ALU_OUT_25_port, DATA_IN(24) => 
                           current_ALU_OUT_24_port, DATA_IN(23) => 
                           current_ALU_OUT_23_port, DATA_IN(22) => 
                           current_ALU_OUT_22_port, DATA_IN(21) => 
                           current_ALU_OUT_21_port, DATA_IN(20) => 
                           current_ALU_OUT_20_port, DATA_IN(19) => 
                           current_ALU_OUT_19_port, DATA_IN(18) => 
                           current_ALU_OUT_18_port, DATA_IN(17) => 
                           current_ALU_OUT_17_port, DATA_IN(16) => 
                           current_ALU_OUT_16_port, DATA_IN(15) => 
                           current_ALU_OUT_15_port, DATA_IN(14) => 
                           current_ALU_OUT_14_port, DATA_IN(13) => 
                           current_ALU_OUT_13_port, DATA_IN(12) => 
                           current_ALU_OUT_12_port, DATA_IN(11) => 
                           current_ALU_OUT_11_port, DATA_IN(10) => 
                           current_ALU_OUT_10_port, DATA_IN(9) => 
                           current_ALU_OUT_9_port, DATA_IN(8) => 
                           current_ALU_OUT_8_port, DATA_IN(7) => 
                           current_ALU_OUT_7_port, DATA_IN(6) => 
                           current_ALU_OUT_6_port, DATA_IN(5) => D_ADDR_5_port,
                           DATA_IN(4) => D_ADDR_4_port, DATA_IN(3) => 
                           D_ADDR_3_port, DATA_IN(2) => D_ADDR_2_port, 
                           DATA_IN(1) => D_ADDR_1_port, DATA_IN(0) => 
                           D_ADDR_0_port, DATA_OUT(31) => 
                           current_ALU_OUT2_31_port, DATA_OUT(30) => 
                           current_ALU_OUT2_30_port, DATA_OUT(29) => 
                           current_ALU_OUT2_29_port, DATA_OUT(28) => 
                           current_ALU_OUT2_28_port, DATA_OUT(27) => 
                           current_ALU_OUT2_27_port, DATA_OUT(26) => 
                           current_ALU_OUT2_26_port, DATA_OUT(25) => 
                           current_ALU_OUT2_25_port, DATA_OUT(24) => 
                           current_ALU_OUT2_24_port, DATA_OUT(23) => 
                           current_ALU_OUT2_23_port, DATA_OUT(22) => 
                           current_ALU_OUT2_22_port, DATA_OUT(21) => 
                           current_ALU_OUT2_21_port, DATA_OUT(20) => 
                           current_ALU_OUT2_20_port, DATA_OUT(19) => 
                           current_ALU_OUT2_19_port, DATA_OUT(18) => 
                           current_ALU_OUT2_18_port, DATA_OUT(17) => 
                           current_ALU_OUT2_17_port, DATA_OUT(16) => 
                           current_ALU_OUT2_16_port, DATA_OUT(15) => 
                           current_ALU_OUT2_15_port, DATA_OUT(14) => 
                           current_ALU_OUT2_14_port, DATA_OUT(13) => 
                           current_ALU_OUT2_13_port, DATA_OUT(12) => 
                           current_ALU_OUT2_12_port, DATA_OUT(11) => 
                           current_ALU_OUT2_11_port, DATA_OUT(10) => 
                           current_ALU_OUT2_10_port, DATA_OUT(9) => 
                           current_ALU_OUT2_9_port, DATA_OUT(8) => 
                           current_ALU_OUT2_8_port, DATA_OUT(7) => 
                           current_ALU_OUT2_7_port, DATA_OUT(6) => 
                           current_ALU_OUT2_6_port, DATA_OUT(5) => 
                           current_ALU_OUT2_5_port, DATA_OUT(4) => 
                           current_ALU_OUT2_4_port, DATA_OUT(3) => 
                           current_ALU_OUT2_3_port, DATA_OUT(2) => 
                           current_ALU_OUT2_2_port, DATA_OUT(1) => 
                           current_ALU_OUT2_1_port, DATA_OUT(0) => 
                           current_ALU_OUT2_0_port);
   BU : BRANCHING_UNIT_N32 port map( CLK => CLK, RST => RST, Reg_A(31) => 
                           A_OUT_31_port, Reg_A(30) => A_OUT_30_port, Reg_A(29)
                           => A_OUT_29_port, Reg_A(28) => A_OUT_28_port, 
                           Reg_A(27) => A_OUT_27_port, Reg_A(26) => 
                           A_OUT_26_port, Reg_A(25) => A_OUT_25_port, Reg_A(24)
                           => A_OUT_24_port, Reg_A(23) => A_OUT_23_port, 
                           Reg_A(22) => A_OUT_22_port, Reg_A(21) => 
                           A_OUT_21_port, Reg_A(20) => A_OUT_20_port, Reg_A(19)
                           => A_OUT_19_port, Reg_A(18) => A_OUT_18_port, 
                           Reg_A(17) => A_OUT_17_port, Reg_A(16) => 
                           A_OUT_16_port, Reg_A(15) => A_OUT_15_port, Reg_A(14)
                           => A_OUT_14_port, Reg_A(13) => A_OUT_13_port, 
                           Reg_A(12) => A_OUT_12_port, Reg_A(11) => 
                           A_OUT_11_port, Reg_A(10) => A_OUT_10_port, Reg_A(9) 
                           => A_OUT_9_port, Reg_A(8) => A_OUT_8_port, Reg_A(7) 
                           => A_OUT_7_port, Reg_A(6) => A_OUT_6_port, Reg_A(5) 
                           => A_OUT_5_port, Reg_A(4) => A_OUT_4_port, Reg_A(3) 
                           => A_OUT_3_port, Reg_A(2) => A_OUT_2_port, Reg_A(1) 
                           => A_OUT_1_port, Reg_A(0) => A_OUT_0_port, EQ_cond 
                           => EQ_COND, IS_JUMP => IS_JUMP, branch_taken => 
                           branch_taken);
   PC_MUX : MUX21_GENERIC_NBIT32_0 port map( A(31) => current_NPC_31_port, 
                           A(30) => current_NPC_30_port, A(29) => 
                           current_NPC_29_port, A(28) => current_NPC_28_port, 
                           A(27) => current_NPC_27_port, A(26) => 
                           current_NPC_26_port, A(25) => current_NPC_25_port, 
                           A(24) => current_NPC_24_port, A(23) => 
                           current_NPC_23_port, A(22) => current_NPC_22_port, 
                           A(21) => current_NPC_21_port, A(20) => 
                           current_NPC_20_port, A(19) => current_NPC_19_port, 
                           A(18) => current_NPC_18_port, A(17) => 
                           current_NPC_17_port, A(16) => current_NPC_16_port, 
                           A(15) => current_NPC_15_port, A(14) => 
                           current_NPC_14_port, A(13) => current_NPC_13_port, 
                           A(12) => current_NPC_12_port, A(11) => 
                           current_NPC_11_port, A(10) => current_NPC_10_port, 
                           A(9) => current_NPC_9_port, A(8) => 
                           current_NPC_8_port, A(7) => current_NPC_7_port, A(6)
                           => current_NPC_6_port, A(5) => current_NPC_5_port, 
                           A(4) => current_NPC_4_port, A(3) => 
                           current_NPC_3_port, A(2) => current_NPC_2_port, A(1)
                           => current_NPC_1_port, A(0) => current_NPC_0_port, 
                           B(31) => current_ALU_OUT_31_port, B(30) => 
                           current_ALU_OUT_30_port, B(29) => 
                           current_ALU_OUT_29_port, B(28) => 
                           current_ALU_OUT_28_port, B(27) => 
                           current_ALU_OUT_27_port, B(26) => 
                           current_ALU_OUT_26_port, B(25) => 
                           current_ALU_OUT_25_port, B(24) => 
                           current_ALU_OUT_24_port, B(23) => 
                           current_ALU_OUT_23_port, B(22) => 
                           current_ALU_OUT_22_port, B(21) => 
                           current_ALU_OUT_21_port, B(20) => 
                           current_ALU_OUT_20_port, B(19) => 
                           current_ALU_OUT_19_port, B(18) => 
                           current_ALU_OUT_18_port, B(17) => 
                           current_ALU_OUT_17_port, B(16) => 
                           current_ALU_OUT_16_port, B(15) => 
                           current_ALU_OUT_15_port, B(14) => 
                           current_ALU_OUT_14_port, B(13) => 
                           current_ALU_OUT_13_port, B(12) => 
                           current_ALU_OUT_12_port, B(11) => 
                           current_ALU_OUT_11_port, B(10) => 
                           current_ALU_OUT_10_port, B(9) => 
                           current_ALU_OUT_9_port, B(8) => 
                           current_ALU_OUT_8_port, B(7) => 
                           current_ALU_OUT_7_port, B(6) => 
                           current_ALU_OUT_6_port, B(5) => D_ADDR_5_port, B(4) 
                           => D_ADDR_4_port, B(3) => D_ADDR_3_port, B(2) => 
                           D_ADDR_2_port, B(1) => D_ADDR_1_port, B(0) => 
                           D_ADDR_0_port, SEL => PC_MUX_SEL, Y(31) => 
                           PC_BUS_31_port, Y(30) => PC_BUS_30_port, Y(29) => 
                           PC_BUS_29_port, Y(28) => PC_BUS_28_port, Y(27) => 
                           PC_BUS_27_port, Y(26) => PC_BUS_26_port, Y(25) => 
                           PC_BUS_25_port, Y(24) => PC_BUS_24_port, Y(23) => 
                           PC_BUS_23_port, Y(22) => PC_BUS_22_port, Y(21) => 
                           PC_BUS_21_port, Y(20) => PC_BUS_20_port, Y(19) => 
                           PC_BUS_19_port, Y(18) => PC_BUS_18_port, Y(17) => 
                           PC_BUS_17_port, Y(16) => PC_BUS_16_port, Y(15) => 
                           PC_BUS_15_port, Y(14) => PC_BUS_14_port, Y(13) => 
                           PC_BUS_13_port, Y(12) => PC_BUS_12_port, Y(11) => 
                           PC_BUS_11_port, Y(10) => PC_BUS_10_port, Y(9) => 
                           PC_BUS_9_port, Y(8) => PC_BUS_8_port, Y(7) => 
                           PC_BUS_7_port, Y(6) => PC_BUS_6_port, Y(5) => 
                           PC_BUS_5_port, Y(4) => PC_BUS_4_port, Y(3) => 
                           PC_BUS_3_port, Y(2) => PC_BUS_2_port, Y(1) => 
                           PC_BUS_1_port, Y(0) => PC_BUS_0_port);
   J_MUX : MUX21 port map( A => X_Logic0_port, B => branch_taken, SEL => 
                           JUMP_EN, Y => PC_MUX_SEL);
   RD_MUX : MUX21_GENERIC_NBIT5_0 port map( A(4) => current_IW_15_port, A(3) =>
                           current_IW_14_port, A(2) => current_IW_13_port, A(1)
                           => current_IW_12_port, A(0) => current_IW_11_port, 
                           B(4) => current_IW_20_port, B(3) => 
                           current_IW_19_port, B(2) => current_IW_18_port, B(1)
                           => current_IW_17_port, B(0) => current_IW_16_port, 
                           SEL => RegIMM_LATCH_EN, Y(4) => WB1_IN_4_port, Y(3) 
                           => WB1_IN_3_port, Y(2) => WB1_IN_2_port, Y(1) => 
                           WB1_IN_1_port, Y(0) => WB1_IN_0_port);
   OP1_MUX : MUX21_GENERIC_NBIT32_4 port map( A(31) => A_OUT_31_port, A(30) => 
                           A_OUT_30_port, A(29) => A_OUT_29_port, A(28) => 
                           A_OUT_28_port, A(27) => A_OUT_27_port, A(26) => 
                           A_OUT_26_port, A(25) => A_OUT_25_port, A(24) => 
                           A_OUT_24_port, A(23) => A_OUT_23_port, A(22) => 
                           A_OUT_22_port, A(21) => A_OUT_21_port, A(20) => 
                           A_OUT_20_port, A(19) => A_OUT_19_port, A(18) => 
                           A_OUT_18_port, A(17) => A_OUT_17_port, A(16) => 
                           A_OUT_16_port, A(15) => A_OUT_15_port, A(14) => 
                           A_OUT_14_port, A(13) => A_OUT_13_port, A(12) => 
                           A_OUT_12_port, A(11) => A_OUT_11_port, A(10) => 
                           A_OUT_10_port, A(9) => A_OUT_9_port, A(8) => 
                           A_OUT_8_port, A(7) => A_OUT_7_port, A(6) => 
                           A_OUT_6_port, A(5) => A_OUT_5_port, A(4) => 
                           A_OUT_4_port, A(3) => A_OUT_3_port, A(2) => 
                           A_OUT_2_port, A(1) => A_OUT_1_port, A(0) => 
                           A_OUT_0_port, B(31) => current_PC1_31_port, B(30) =>
                           current_PC1_30_port, B(29) => current_PC1_29_port, 
                           B(28) => current_PC1_28_port, B(27) => 
                           current_PC1_27_port, B(26) => current_PC1_26_port, 
                           B(25) => current_PC1_25_port, B(24) => 
                           current_PC1_24_port, B(23) => current_PC1_23_port, 
                           B(22) => current_PC1_22_port, B(21) => 
                           current_PC1_21_port, B(20) => current_PC1_20_port, 
                           B(19) => current_PC1_19_port, B(18) => 
                           current_PC1_18_port, B(17) => current_PC1_17_port, 
                           B(16) => current_PC1_16_port, B(15) => 
                           current_PC1_15_port, B(14) => current_PC1_14_port, 
                           B(13) => current_PC1_13_port, B(12) => 
                           current_PC1_12_port, B(11) => current_PC1_11_port, 
                           B(10) => current_PC1_10_port, B(9) => 
                           current_PC1_9_port, B(8) => current_PC1_8_port, B(7)
                           => current_PC1_7_port, B(6) => current_PC1_6_port, 
                           B(5) => current_PC1_5_port, B(4) => 
                           current_PC1_4_port, B(3) => current_PC1_3_port, B(2)
                           => current_PC1_2_port, B(1) => current_PC1_1_port, 
                           B(0) => current_PC1_0_port, SEL => MUXA_SEL, Y(31) 
                           => ALU_OP1_31_port, Y(30) => ALU_OP1_30_port, Y(29) 
                           => ALU_OP1_29_port, Y(28) => ALU_OP1_28_port, Y(27) 
                           => ALU_OP1_27_port, Y(26) => ALU_OP1_26_port, Y(25) 
                           => ALU_OP1_25_port, Y(24) => ALU_OP1_24_port, Y(23) 
                           => ALU_OP1_23_port, Y(22) => ALU_OP1_22_port, Y(21) 
                           => ALU_OP1_21_port, Y(20) => ALU_OP1_20_port, Y(19) 
                           => ALU_OP1_19_port, Y(18) => ALU_OP1_18_port, Y(17) 
                           => ALU_OP1_17_port, Y(16) => ALU_OP1_16_port, Y(15) 
                           => ALU_OP1_15_port, Y(14) => ALU_OP1_14_port, Y(13) 
                           => ALU_OP1_13_port, Y(12) => ALU_OP1_12_port, Y(11) 
                           => ALU_OP1_11_port, Y(10) => ALU_OP1_10_port, Y(9) 
                           => ALU_OP1_9_port, Y(8) => ALU_OP1_8_port, Y(7) => 
                           ALU_OP1_7_port, Y(6) => ALU_OP1_6_port, Y(5) => 
                           ALU_OP1_5_port, Y(4) => ALU_OP1_4_port, Y(3) => 
                           ALU_OP1_3_port, Y(2) => ALU_OP1_2_port, Y(1) => 
                           ALU_OP1_1_port, Y(0) => ALU_OP1_0_port);
   OP2_MUX : MUX21_GENERIC_NBIT32_3 port map( A(31) => B_OUT_31_port, A(30) => 
                           B_OUT_30_port, A(29) => B_OUT_29_port, A(28) => 
                           B_OUT_28_port, A(27) => B_OUT_27_port, A(26) => 
                           B_OUT_26_port, A(25) => B_OUT_25_port, A(24) => 
                           B_OUT_24_port, A(23) => B_OUT_23_port, A(22) => 
                           B_OUT_22_port, A(21) => B_OUT_21_port, A(20) => 
                           B_OUT_20_port, A(19) => B_OUT_19_port, A(18) => 
                           B_OUT_18_port, A(17) => B_OUT_17_port, A(16) => 
                           B_OUT_16_port, A(15) => B_OUT_15_port, A(14) => 
                           B_OUT_14_port, A(13) => B_OUT_13_port, A(12) => 
                           B_OUT_12_port, A(11) => B_OUT_11_port, A(10) => 
                           B_OUT_10_port, A(9) => B_OUT_9_port, A(8) => 
                           B_OUT_8_port, A(7) => B_OUT_7_port, A(6) => 
                           B_OUT_6_port, A(5) => B_OUT_5_port, A(4) => 
                           B_OUT_4_port, A(3) => B_OUT_3_port, A(2) => 
                           B_OUT_2_port, A(1) => B_OUT_1_port, A(0) => 
                           B_OUT_0_port, B(31) => IMM_OUT_31_port, B(30) => 
                           IMM_OUT_30_port, B(29) => IMM_OUT_29_port, B(28) => 
                           IMM_OUT_28_port, B(27) => IMM_OUT_27_port, B(26) => 
                           IMM_OUT_26_port, B(25) => IMM_OUT_25_port, B(24) => 
                           IMM_OUT_24_port, B(23) => IMM_OUT_23_port, B(22) => 
                           IMM_OUT_22_port, B(21) => IMM_OUT_21_port, B(20) => 
                           IMM_OUT_20_port, B(19) => IMM_OUT_19_port, B(18) => 
                           IMM_OUT_18_port, B(17) => IMM_OUT_17_port, B(16) => 
                           IMM_OUT_16_port, B(15) => IMM_OUT_15_port, B(14) => 
                           IMM_OUT_14_port, B(13) => IMM_OUT_13_port, B(12) => 
                           IMM_OUT_12_port, B(11) => IMM_OUT_11_port, B(10) => 
                           IMM_OUT_10_port, B(9) => IMM_OUT_9_port, B(8) => 
                           IMM_OUT_8_port, B(7) => IMM_OUT_7_port, B(6) => 
                           IMM_OUT_6_port, B(5) => IMM_OUT_5_port, B(4) => 
                           IMM_OUT_4_port, B(3) => IMM_OUT_3_port, B(2) => 
                           IMM_OUT_2_port, B(1) => IMM_OUT_1_port, B(0) => 
                           IMM_OUT_0_port, SEL => MUXB_SEL, Y(31) => 
                           ALU_OP2_31_port, Y(30) => ALU_OP2_30_port, Y(29) => 
                           ALU_OP2_29_port, Y(28) => ALU_OP2_28_port, Y(27) => 
                           ALU_OP2_27_port, Y(26) => ALU_OP2_26_port, Y(25) => 
                           ALU_OP2_25_port, Y(24) => ALU_OP2_24_port, Y(23) => 
                           ALU_OP2_23_port, Y(22) => ALU_OP2_22_port, Y(21) => 
                           ALU_OP2_21_port, Y(20) => ALU_OP2_20_port, Y(19) => 
                           ALU_OP2_19_port, Y(18) => ALU_OP2_18_port, Y(17) => 
                           ALU_OP2_17_port, Y(16) => ALU_OP2_16_port, Y(15) => 
                           ALU_OP2_15_port, Y(14) => ALU_OP2_14_port, Y(13) => 
                           ALU_OP2_13_port, Y(12) => ALU_OP2_12_port, Y(11) => 
                           ALU_OP2_11_port, Y(10) => ALU_OP2_10_port, Y(9) => 
                           ALU_OP2_9_port, Y(8) => ALU_OP2_8_port, Y(7) => 
                           ALU_OP2_7_port, Y(6) => ALU_OP2_6_port, Y(5) => 
                           ALU_OP2_5_port, Y(4) => ALU_OP2_4_port, Y(3) => 
                           ALU_OP2_3_port, Y(2) => ALU_OP2_2_port, Y(1) => 
                           ALU_OP2_1_port, Y(0) => ALU_OP2_0_port);
   OUT_MUX : MUX21_GENERIC_NBIT32_2 port map( A(31) => D_DATA_OUT(31), A(30) =>
                           D_DATA_OUT(30), A(29) => D_DATA_OUT(29), A(28) => 
                           D_DATA_OUT(28), A(27) => D_DATA_OUT(27), A(26) => 
                           D_DATA_OUT(26), A(25) => D_DATA_OUT(25), A(24) => 
                           D_DATA_OUT(24), A(23) => D_DATA_OUT(23), A(22) => 
                           D_DATA_OUT(22), A(21) => D_DATA_OUT(21), A(20) => 
                           D_DATA_OUT(20), A(19) => D_DATA_OUT(19), A(18) => 
                           D_DATA_OUT(18), A(17) => D_DATA_OUT(17), A(16) => 
                           D_DATA_OUT(16), A(15) => D_DATA_OUT(15), A(14) => 
                           D_DATA_OUT(14), A(13) => D_DATA_OUT(13), A(12) => 
                           D_DATA_OUT(12), A(11) => D_DATA_OUT(11), A(10) => 
                           D_DATA_OUT(10), A(9) => D_DATA_OUT(9), A(8) => 
                           D_DATA_OUT(8), A(7) => D_DATA_OUT(7), A(6) => 
                           D_DATA_OUT(6), A(5) => D_DATA_OUT(5), A(4) => 
                           D_DATA_OUT(4), A(3) => D_DATA_OUT(3), A(2) => 
                           D_DATA_OUT(2), A(1) => D_DATA_OUT(1), A(0) => 
                           D_DATA_OUT(0), B(31) => current_ALU_OUT2_31_port, 
                           B(30) => current_ALU_OUT2_30_port, B(29) => 
                           current_ALU_OUT2_29_port, B(28) => 
                           current_ALU_OUT2_28_port, B(27) => 
                           current_ALU_OUT2_27_port, B(26) => 
                           current_ALU_OUT2_26_port, B(25) => 
                           current_ALU_OUT2_25_port, B(24) => 
                           current_ALU_OUT2_24_port, B(23) => 
                           current_ALU_OUT2_23_port, B(22) => 
                           current_ALU_OUT2_22_port, B(21) => 
                           current_ALU_OUT2_21_port, B(20) => 
                           current_ALU_OUT2_20_port, B(19) => 
                           current_ALU_OUT2_19_port, B(18) => 
                           current_ALU_OUT2_18_port, B(17) => 
                           current_ALU_OUT2_17_port, B(16) => 
                           current_ALU_OUT2_16_port, B(15) => 
                           current_ALU_OUT2_15_port, B(14) => 
                           current_ALU_OUT2_14_port, B(13) => 
                           current_ALU_OUT2_13_port, B(12) => 
                           current_ALU_OUT2_12_port, B(11) => 
                           current_ALU_OUT2_11_port, B(10) => 
                           current_ALU_OUT2_10_port, B(9) => 
                           current_ALU_OUT2_9_port, B(8) => 
                           current_ALU_OUT2_8_port, B(7) => 
                           current_ALU_OUT2_7_port, B(6) => 
                           current_ALU_OUT2_6_port, B(5) => 
                           current_ALU_OUT2_5_port, B(4) => 
                           current_ALU_OUT2_4_port, B(3) => 
                           current_ALU_OUT2_3_port, B(2) => 
                           current_ALU_OUT2_2_port, B(1) => 
                           current_ALU_OUT2_1_port, B(0) => 
                           current_ALU_OUT2_0_port, SEL => WB_MUX_SEL, Y(31) =>
                           OUT_MUX_DATA_31_port, Y(30) => OUT_MUX_DATA_30_port,
                           Y(29) => OUT_MUX_DATA_29_port, Y(28) => 
                           OUT_MUX_DATA_28_port, Y(27) => OUT_MUX_DATA_27_port,
                           Y(26) => OUT_MUX_DATA_26_port, Y(25) => 
                           OUT_MUX_DATA_25_port, Y(24) => OUT_MUX_DATA_24_port,
                           Y(23) => OUT_MUX_DATA_23_port, Y(22) => 
                           OUT_MUX_DATA_22_port, Y(21) => OUT_MUX_DATA_21_port,
                           Y(20) => OUT_MUX_DATA_20_port, Y(19) => 
                           OUT_MUX_DATA_19_port, Y(18) => OUT_MUX_DATA_18_port,
                           Y(17) => OUT_MUX_DATA_17_port, Y(16) => 
                           OUT_MUX_DATA_16_port, Y(15) => OUT_MUX_DATA_15_port,
                           Y(14) => OUT_MUX_DATA_14_port, Y(13) => 
                           OUT_MUX_DATA_13_port, Y(12) => OUT_MUX_DATA_12_port,
                           Y(11) => OUT_MUX_DATA_11_port, Y(10) => 
                           OUT_MUX_DATA_10_port, Y(9) => OUT_MUX_DATA_9_port, 
                           Y(8) => OUT_MUX_DATA_8_port, Y(7) => 
                           OUT_MUX_DATA_7_port, Y(6) => OUT_MUX_DATA_6_port, 
                           Y(5) => OUT_MUX_DATA_5_port, Y(4) => 
                           OUT_MUX_DATA_4_port, Y(3) => OUT_MUX_DATA_3_port, 
                           Y(2) => OUT_MUX_DATA_2_port, Y(1) => 
                           OUT_MUX_DATA_1_port, Y(0) => OUT_MUX_DATA_0_port);
   JAL_DATA_MUX : MUX21_GENERIC_NBIT32_1 port map( A(31) => 
                           OUT_MUX_DATA_31_port, A(30) => OUT_MUX_DATA_30_port,
                           A(29) => OUT_MUX_DATA_29_port, A(28) => 
                           OUT_MUX_DATA_28_port, A(27) => OUT_MUX_DATA_27_port,
                           A(26) => OUT_MUX_DATA_26_port, A(25) => 
                           OUT_MUX_DATA_25_port, A(24) => OUT_MUX_DATA_24_port,
                           A(23) => OUT_MUX_DATA_23_port, A(22) => 
                           OUT_MUX_DATA_22_port, A(21) => OUT_MUX_DATA_21_port,
                           A(20) => OUT_MUX_DATA_20_port, A(19) => 
                           OUT_MUX_DATA_19_port, A(18) => OUT_MUX_DATA_18_port,
                           A(17) => OUT_MUX_DATA_17_port, A(16) => 
                           OUT_MUX_DATA_16_port, A(15) => OUT_MUX_DATA_15_port,
                           A(14) => OUT_MUX_DATA_14_port, A(13) => 
                           OUT_MUX_DATA_13_port, A(12) => OUT_MUX_DATA_12_port,
                           A(11) => OUT_MUX_DATA_11_port, A(10) => 
                           OUT_MUX_DATA_10_port, A(9) => OUT_MUX_DATA_9_port, 
                           A(8) => OUT_MUX_DATA_8_port, A(7) => 
                           OUT_MUX_DATA_7_port, A(6) => OUT_MUX_DATA_6_port, 
                           A(5) => OUT_MUX_DATA_5_port, A(4) => 
                           OUT_MUX_DATA_4_port, A(3) => OUT_MUX_DATA_3_port, 
                           A(2) => OUT_MUX_DATA_2_port, A(1) => 
                           OUT_MUX_DATA_1_port, A(0) => OUT_MUX_DATA_0_port, 
                           B(31) => current_PC3_31_port, B(30) => 
                           current_PC3_30_port, B(29) => current_PC3_29_port, 
                           B(28) => current_PC3_28_port, B(27) => 
                           current_PC3_27_port, B(26) => current_PC3_26_port, 
                           B(25) => current_PC3_25_port, B(24) => 
                           current_PC3_24_port, B(23) => current_PC3_23_port, 
                           B(22) => current_PC3_22_port, B(21) => 
                           current_PC3_21_port, B(20) => current_PC3_20_port, 
                           B(19) => current_PC3_19_port, B(18) => 
                           current_PC3_18_port, B(17) => current_PC3_17_port, 
                           B(16) => current_PC3_16_port, B(15) => 
                           current_PC3_15_port, B(14) => current_PC3_14_port, 
                           B(13) => current_PC3_13_port, B(12) => 
                           current_PC3_12_port, B(11) => current_PC3_11_port, 
                           B(10) => current_PC3_10_port, B(9) => 
                           current_PC3_9_port, B(8) => current_PC3_8_port, B(7)
                           => current_PC3_7_port, B(6) => current_PC3_6_port, 
                           B(5) => current_PC3_5_port, B(4) => 
                           current_PC3_4_port, B(3) => current_PC3_3_port, B(2)
                           => current_PC3_2_port, B(1) => current_PC3_1_port, 
                           B(0) => current_PC3_0_port, SEL => IS_JAL, Y(31) => 
                           WB_DATA_31_port, Y(30) => WB_DATA_30_port, Y(29) => 
                           WB_DATA_29_port, Y(28) => WB_DATA_28_port, Y(27) => 
                           WB_DATA_27_port, Y(26) => WB_DATA_26_port, Y(25) => 
                           WB_DATA_25_port, Y(24) => WB_DATA_24_port, Y(23) => 
                           WB_DATA_23_port, Y(22) => WB_DATA_22_port, Y(21) => 
                           WB_DATA_21_port, Y(20) => WB_DATA_20_port, Y(19) => 
                           WB_DATA_19_port, Y(18) => WB_DATA_18_port, Y(17) => 
                           WB_DATA_17_port, Y(16) => WB_DATA_16_port, Y(15) => 
                           WB_DATA_15_port, Y(14) => WB_DATA_14_port, Y(13) => 
                           WB_DATA_13_port, Y(12) => WB_DATA_12_port, Y(11) => 
                           WB_DATA_11_port, Y(10) => WB_DATA_10_port, Y(9) => 
                           WB_DATA_9_port, Y(8) => WB_DATA_8_port, Y(7) => 
                           WB_DATA_7_port, Y(6) => WB_DATA_6_port, Y(5) => 
                           WB_DATA_5_port, Y(4) => WB_DATA_4_port, Y(3) => 
                           WB_DATA_3_port, Y(2) => WB_DATA_2_port, Y(1) => 
                           WB_DATA_1_port, Y(0) => WB_DATA_0_port);
   JAL_ADDR_MUX : MUX21_GENERIC_NBIT5_1 port map( A(4) => WB3_OUT_4_port, A(3) 
                           => WB3_OUT_3_port, A(2) => WB3_OUT_2_port, A(1) => 
                           WB3_OUT_1_port, A(0) => WB3_OUT_0_port, B(4) => 
                           X_Logic1_port, B(3) => X_Logic1_port, B(2) => 
                           X_Logic1_port, B(1) => X_Logic1_port, B(0) => 
                           X_Logic1_port, SEL => IS_JAL, Y(4) => WB_ADDR_4_port
                           , Y(3) => WB_ADDR_3_port, Y(2) => WB_ADDR_2_port, 
                           Y(1) => WB_ADDR_1_port, Y(0) => WB_ADDR_0_port);
   PC_ADDER : ADDER_N32 port map( CURR_ADDR(31) => current_PC_31_port, 
                           CURR_ADDR(30) => current_PC_30_port, CURR_ADDR(29) 
                           => current_PC_29_port, CURR_ADDR(28) => 
                           current_PC_28_port, CURR_ADDR(27) => 
                           current_PC_27_port, CURR_ADDR(26) => 
                           current_PC_26_port, CURR_ADDR(25) => 
                           current_PC_25_port, CURR_ADDR(24) => 
                           current_PC_24_port, CURR_ADDR(23) => 
                           current_PC_23_port, CURR_ADDR(22) => 
                           current_PC_22_port, CURR_ADDR(21) => 
                           current_PC_21_port, CURR_ADDR(20) => 
                           current_PC_20_port, CURR_ADDR(19) => 
                           current_PC_19_port, CURR_ADDR(18) => 
                           current_PC_18_port, CURR_ADDR(17) => 
                           current_PC_17_port, CURR_ADDR(16) => 
                           current_PC_16_port, CURR_ADDR(15) => 
                           current_PC_15_port, CURR_ADDR(14) => 
                           current_PC_14_port, CURR_ADDR(13) => 
                           current_PC_13_port, CURR_ADDR(12) => 
                           current_PC_12_port, CURR_ADDR(11) => 
                           current_PC_11_port, CURR_ADDR(10) => 
                           current_PC_10_port, CURR_ADDR(9) => 
                           current_PC_9_port, CURR_ADDR(8) => current_PC_8_port
                           , CURR_ADDR(7) => current_PC_7_port, CURR_ADDR(6) =>
                           current_PC_6_port, CURR_ADDR(5) => current_PC_5_port
                           , CURR_ADDR(4) => current_PC_4_port, CURR_ADDR(3) =>
                           current_PC_3_port, CURR_ADDR(2) => current_PC_2_port
                           , CURR_ADDR(1) => current_PC_1_port, CURR_ADDR(0) =>
                           current_PC_0_port, NEXT_ADDR(31) => next_NPC_31_port
                           , NEXT_ADDR(30) => next_NPC_30_port, NEXT_ADDR(29) 
                           => next_NPC_29_port, NEXT_ADDR(28) => 
                           next_NPC_28_port, NEXT_ADDR(27) => next_NPC_27_port,
                           NEXT_ADDR(26) => next_NPC_26_port, NEXT_ADDR(25) => 
                           next_NPC_25_port, NEXT_ADDR(24) => next_NPC_24_port,
                           NEXT_ADDR(23) => next_NPC_23_port, NEXT_ADDR(22) => 
                           next_NPC_22_port, NEXT_ADDR(21) => next_NPC_21_port,
                           NEXT_ADDR(20) => next_NPC_20_port, NEXT_ADDR(19) => 
                           next_NPC_19_port, NEXT_ADDR(18) => next_NPC_18_port,
                           NEXT_ADDR(17) => next_NPC_17_port, NEXT_ADDR(16) => 
                           next_NPC_16_port, NEXT_ADDR(15) => next_NPC_15_port,
                           NEXT_ADDR(14) => next_NPC_14_port, NEXT_ADDR(13) => 
                           next_NPC_13_port, NEXT_ADDR(12) => next_NPC_12_port,
                           NEXT_ADDR(11) => next_NPC_11_port, NEXT_ADDR(10) => 
                           next_NPC_10_port, NEXT_ADDR(9) => next_NPC_9_port, 
                           NEXT_ADDR(8) => next_NPC_8_port, NEXT_ADDR(7) => 
                           next_NPC_7_port, NEXT_ADDR(6) => next_NPC_6_port, 
                           NEXT_ADDR(5) => next_NPC_5_port, NEXT_ADDR(4) => 
                           next_NPC_4_port, NEXT_ADDR(3) => next_NPC_3_port, 
                           NEXT_ADDR(2) => next_NPC_2_port, NEXT_ADDR(1) => 
                           next_NPC_1_port, NEXT_ADDR(0) => next_NPC_0_port);
   EXT : EXTENDER_NBIT32_IMM_field_lenght16 port map( NOT_EXT_IMM(15) => 
                           IMM_IN_15_port, NOT_EXT_IMM(14) => IMM_IN_14_port, 
                           NOT_EXT_IMM(13) => IMM_IN_13_port, NOT_EXT_IMM(12) 
                           => IMM_IN_12_port, NOT_EXT_IMM(11) => IMM_IN_11_port
                           , NOT_EXT_IMM(10) => IMM_IN_10_port, NOT_EXT_IMM(9) 
                           => IMM_IN_9_port, NOT_EXT_IMM(8) => IMM_IN_8_port, 
                           NOT_EXT_IMM(7) => IMM_IN_7_port, NOT_EXT_IMM(6) => 
                           IMM_IN_6_port, NOT_EXT_IMM(5) => IMM_IN_5_port, 
                           NOT_EXT_IMM(4) => IMM_IN_4_port, NOT_EXT_IMM(3) => 
                           IMM_IN_3_port, NOT_EXT_IMM(2) => IMM_IN_2_port, 
                           NOT_EXT_IMM(1) => IMM_IN_1_port, NOT_EXT_IMM(0) => 
                           IMM_IN_0_port, SIGNED_IMM => SIGNED_IMM, EXT_IMM(31)
                           => IMM_OUT_31_port, EXT_IMM(30) => IMM_OUT_30_port, 
                           EXT_IMM(29) => IMM_OUT_29_port, EXT_IMM(28) => 
                           IMM_OUT_28_port, EXT_IMM(27) => IMM_OUT_27_port, 
                           EXT_IMM(26) => IMM_OUT_26_port, EXT_IMM(25) => 
                           IMM_OUT_25_port, EXT_IMM(24) => IMM_OUT_24_port, 
                           EXT_IMM(23) => IMM_OUT_23_port, EXT_IMM(22) => 
                           IMM_OUT_22_port, EXT_IMM(21) => IMM_OUT_21_port, 
                           EXT_IMM(20) => IMM_OUT_20_port, EXT_IMM(19) => 
                           IMM_OUT_19_port, EXT_IMM(18) => IMM_OUT_18_port, 
                           EXT_IMM(17) => IMM_OUT_17_port, EXT_IMM(16) => 
                           IMM_OUT_16_port, EXT_IMM(15) => IMM_OUT_15_port, 
                           EXT_IMM(14) => IMM_OUT_14_port, EXT_IMM(13) => 
                           IMM_OUT_13_port, EXT_IMM(12) => IMM_OUT_12_port, 
                           EXT_IMM(11) => IMM_OUT_11_port, EXT_IMM(10) => 
                           IMM_OUT_10_port, EXT_IMM(9) => IMM_OUT_9_port, 
                           EXT_IMM(8) => IMM_OUT_8_port, EXT_IMM(7) => 
                           IMM_OUT_7_port, EXT_IMM(6) => IMM_OUT_6_port, 
                           EXT_IMM(5) => IMM_OUT_5_port, EXT_IMM(4) => 
                           IMM_OUT_4_port, EXT_IMM(3) => IMM_OUT_3_port, 
                           EXT_IMM(2) => IMM_OUT_2_port, EXT_IMM(1) => 
                           IMM_OUT_1_port, EXT_IMM(0) => IMM_OUT_0_port);
   ALU_i : ALU_N32 port map( FUNC(0) => ALU_OPCODE(0), FUNC(1) => ALU_OPCODE(1)
                           , FUNC(2) => ALU_OPCODE(2), FUNC(3) => ALU_OPCODE(3)
                           , DATA1(31) => ALU_OP1_31_port, DATA1(30) => 
                           ALU_OP1_30_port, DATA1(29) => ALU_OP1_29_port, 
                           DATA1(28) => ALU_OP1_28_port, DATA1(27) => 
                           ALU_OP1_27_port, DATA1(26) => ALU_OP1_26_port, 
                           DATA1(25) => ALU_OP1_25_port, DATA1(24) => 
                           ALU_OP1_24_port, DATA1(23) => ALU_OP1_23_port, 
                           DATA1(22) => ALU_OP1_22_port, DATA1(21) => 
                           ALU_OP1_21_port, DATA1(20) => ALU_OP1_20_port, 
                           DATA1(19) => ALU_OP1_19_port, DATA1(18) => 
                           ALU_OP1_18_port, DATA1(17) => ALU_OP1_17_port, 
                           DATA1(16) => ALU_OP1_16_port, DATA1(15) => 
                           ALU_OP1_15_port, DATA1(14) => ALU_OP1_14_port, 
                           DATA1(13) => ALU_OP1_13_port, DATA1(12) => 
                           ALU_OP1_12_port, DATA1(11) => ALU_OP1_11_port, 
                           DATA1(10) => ALU_OP1_10_port, DATA1(9) => 
                           ALU_OP1_9_port, DATA1(8) => ALU_OP1_8_port, DATA1(7)
                           => ALU_OP1_7_port, DATA1(6) => ALU_OP1_6_port, 
                           DATA1(5) => ALU_OP1_5_port, DATA1(4) => 
                           ALU_OP1_4_port, DATA1(3) => ALU_OP1_3_port, DATA1(2)
                           => ALU_OP1_2_port, DATA1(1) => ALU_OP1_1_port, 
                           DATA1(0) => ALU_OP1_0_port, DATA2(31) => 
                           ALU_OP2_31_port, DATA2(30) => ALU_OP2_30_port, 
                           DATA2(29) => ALU_OP2_29_port, DATA2(28) => 
                           ALU_OP2_28_port, DATA2(27) => ALU_OP2_27_port, 
                           DATA2(26) => ALU_OP2_26_port, DATA2(25) => 
                           ALU_OP2_25_port, DATA2(24) => ALU_OP2_24_port, 
                           DATA2(23) => ALU_OP2_23_port, DATA2(22) => 
                           ALU_OP2_22_port, DATA2(21) => ALU_OP2_21_port, 
                           DATA2(20) => ALU_OP2_20_port, DATA2(19) => 
                           ALU_OP2_19_port, DATA2(18) => ALU_OP2_18_port, 
                           DATA2(17) => ALU_OP2_17_port, DATA2(16) => 
                           ALU_OP2_16_port, DATA2(15) => ALU_OP2_15_port, 
                           DATA2(14) => ALU_OP2_14_port, DATA2(13) => 
                           ALU_OP2_13_port, DATA2(12) => ALU_OP2_12_port, 
                           DATA2(11) => ALU_OP2_11_port, DATA2(10) => 
                           ALU_OP2_10_port, DATA2(9) => ALU_OP2_9_port, 
                           DATA2(8) => ALU_OP2_8_port, DATA2(7) => 
                           ALU_OP2_7_port, DATA2(6) => ALU_OP2_6_port, DATA2(5)
                           => ALU_OP2_5_port, DATA2(4) => ALU_OP2_4_port, 
                           DATA2(3) => ALU_OP2_3_port, DATA2(2) => 
                           ALU_OP2_2_port, DATA2(1) => ALU_OP2_1_port, DATA2(0)
                           => ALU_OP2_0_port, OUTALU(31) => 
                           next_ALU_OUT_31_port, OUTALU(30) => 
                           next_ALU_OUT_30_port, OUTALU(29) => 
                           next_ALU_OUT_29_port, OUTALU(28) => 
                           next_ALU_OUT_28_port, OUTALU(27) => 
                           next_ALU_OUT_27_port, OUTALU(26) => 
                           next_ALU_OUT_26_port, OUTALU(25) => 
                           next_ALU_OUT_25_port, OUTALU(24) => 
                           next_ALU_OUT_24_port, OUTALU(23) => 
                           next_ALU_OUT_23_port, OUTALU(22) => 
                           next_ALU_OUT_22_port, OUTALU(21) => 
                           next_ALU_OUT_21_port, OUTALU(20) => 
                           next_ALU_OUT_20_port, OUTALU(19) => 
                           next_ALU_OUT_19_port, OUTALU(18) => 
                           next_ALU_OUT_18_port, OUTALU(17) => 
                           next_ALU_OUT_17_port, OUTALU(16) => 
                           next_ALU_OUT_16_port, OUTALU(15) => 
                           next_ALU_OUT_15_port, OUTALU(14) => 
                           next_ALU_OUT_14_port, OUTALU(13) => 
                           next_ALU_OUT_13_port, OUTALU(12) => 
                           next_ALU_OUT_12_port, OUTALU(11) => 
                           next_ALU_OUT_11_port, OUTALU(10) => 
                           next_ALU_OUT_10_port, OUTALU(9) => 
                           next_ALU_OUT_9_port, OUTALU(8) => 
                           next_ALU_OUT_8_port, OUTALU(7) => 
                           next_ALU_OUT_7_port, OUTALU(6) => 
                           next_ALU_OUT_6_port, OUTALU(5) => 
                           next_ALU_OUT_5_port, OUTALU(4) => 
                           next_ALU_OUT_4_port, OUTALU(3) => 
                           next_ALU_OUT_3_port, OUTALU(2) => 
                           next_ALU_OUT_2_port, OUTALU(1) => 
                           next_ALU_OUT_1_port, OUTALU(0) => 
                           next_ALU_OUT_0_port);
   U3 : AND2_X1 port map( A1 => PC_LATCH_EN, A2 => PC_BUS_9_port, ZN => 
                           current_PC_9_port);
   U4 : AND2_X1 port map( A1 => PC_BUS_8_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_8_port);
   U5 : AND2_X1 port map( A1 => PC_BUS_7_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_7_port);
   U6 : AND2_X1 port map( A1 => PC_BUS_6_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_6_port);
   U7 : AND2_X1 port map( A1 => PC_BUS_5_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_5_port);
   U8 : AND2_X1 port map( A1 => PC_BUS_4_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_4_port);
   U9 : AND2_X1 port map( A1 => PC_BUS_3_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_3_port);
   U10 : AND2_X1 port map( A1 => PC_BUS_31_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_31_port);
   U11 : AND2_X1 port map( A1 => PC_BUS_30_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_30_port);
   U12 : AND2_X1 port map( A1 => PC_BUS_2_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_2_port);
   U13 : AND2_X1 port map( A1 => PC_BUS_29_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_29_port);
   U14 : AND2_X1 port map( A1 => PC_BUS_28_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_28_port);
   U15 : AND2_X1 port map( A1 => PC_BUS_27_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_27_port);
   U16 : AND2_X1 port map( A1 => PC_BUS_26_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_26_port);
   U17 : AND2_X1 port map( A1 => PC_BUS_25_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_25_port);
   U18 : AND2_X1 port map( A1 => PC_BUS_24_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_24_port);
   U19 : AND2_X1 port map( A1 => PC_BUS_23_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_23_port);
   U20 : AND2_X1 port map( A1 => PC_BUS_22_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_22_port);
   U21 : AND2_X1 port map( A1 => PC_BUS_21_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_21_port);
   U22 : AND2_X1 port map( A1 => PC_BUS_20_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_20_port);
   U23 : AND2_X1 port map( A1 => PC_BUS_1_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_1_port);
   U24 : AND2_X1 port map( A1 => PC_BUS_19_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_19_port);
   U25 : AND2_X1 port map( A1 => PC_BUS_18_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_18_port);
   U26 : AND2_X1 port map( A1 => PC_BUS_17_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_17_port);
   U27 : AND2_X1 port map( A1 => PC_BUS_16_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_16_port);
   U28 : AND2_X1 port map( A1 => PC_BUS_15_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_15_port);
   U29 : AND2_X1 port map( A1 => PC_BUS_14_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_14_port);
   U30 : AND2_X1 port map( A1 => PC_BUS_13_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_13_port);
   U31 : AND2_X1 port map( A1 => PC_BUS_12_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_12_port);
   U32 : AND2_X1 port map( A1 => PC_BUS_11_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_11_port);
   U33 : AND2_X1 port map( A1 => PC_BUS_10_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_10_port);
   U34 : AND2_X1 port map( A1 => PC_BUS_0_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_0_port);

end SYN_STRUCTURE;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_0 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_0;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( CLK, RST : in std_logic;  I_ADDR : out std_logic_vector (31 downto 0);
         I_DATA : in std_logic_vector (31 downto 0);  D_RR, D_WR : out 
         std_logic;  D_ADDR : out std_logic_vector (5 downto 0);  D_DATA_IN : 
         out std_logic_vector (31 downto 0);  D_DATA_OUT : in std_logic_vector 
         (31 downto 0));

end DLX;

architecture SYN_DLX_RTL of DLX is

   component dlx_cu
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
            EQ_COND, IS_JUMP : out std_logic;  ALU_OPCODE : out 
            std_logic_vector (0 to 3);  DRAM_WE, LMD_LATCH_EN, JUMP_EN, 
            PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE : out std_logic);
   end component;
   
   component DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64
      port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
            EQ_COND, IS_JUMP : in std_logic;  ALU_OPCODE : in std_logic_vector 
            (0 to 3);  JUMP_EN, PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE : in 
            std_logic;  D_ADDR : out std_logic_vector (5 downto 0);  D_DATA_IN 
            : out std_logic_vector (31 downto 0);  D_DATA_OUT, PC_IN : in 
            std_logic_vector (31 downto 0);  PC_BUS : out std_logic_vector (31 
            downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_0
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal I_ADDR_31_port, I_ADDR_30_port, I_ADDR_29_port, I_ADDR_28_port, 
      I_ADDR_27_port, I_ADDR_26_port, I_ADDR_25_port, I_ADDR_24_port, 
      I_ADDR_23_port, I_ADDR_22_port, I_ADDR_21_port, I_ADDR_20_port, 
      I_ADDR_19_port, I_ADDR_18_port, I_ADDR_17_port, I_ADDR_16_port, 
      I_ADDR_15_port, I_ADDR_14_port, I_ADDR_13_port, I_ADDR_12_port, 
      I_ADDR_11_port, I_ADDR_10_port, I_ADDR_9_port, I_ADDR_8_port, 
      I_ADDR_7_port, I_ADDR_6_port, I_ADDR_5_port, I_ADDR_4_port, I_ADDR_3_port
      , I_ADDR_2_port, I_ADDR_1_port, I_ADDR_0_port, PC_LATCH_EN, 
      PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, IR_LATCH_EN, NPC_LATCH_EN,
      RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, 
      MUXB_SEL, ALU_OUTREG_EN, EQ_COND, IS_JUMP, ALU_OPCODE_3_port, 
      ALU_OPCODE_2_port, ALU_OPCODE_1_port, ALU_OPCODE_0_port, JUMP_EN, IS_JAL,
      WB_MUX_SEL, RF_WE, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164
      , n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173,
      n_2174, n_2175 : std_logic;

begin
   I_ADDR <= ( I_ADDR_31_port, I_ADDR_30_port, I_ADDR_29_port, I_ADDR_28_port, 
      I_ADDR_27_port, I_ADDR_26_port, I_ADDR_25_port, I_ADDR_24_port, 
      I_ADDR_23_port, I_ADDR_22_port, I_ADDR_21_port, I_ADDR_20_port, 
      I_ADDR_19_port, I_ADDR_18_port, I_ADDR_17_port, I_ADDR_16_port, 
      I_ADDR_15_port, I_ADDR_14_port, I_ADDR_13_port, I_ADDR_12_port, 
      I_ADDR_11_port, I_ADDR_10_port, I_ADDR_9_port, I_ADDR_8_port, 
      I_ADDR_7_port, I_ADDR_6_port, I_ADDR_5_port, I_ADDR_4_port, I_ADDR_3_port
      , I_ADDR_2_port, I_ADDR_1_port, I_ADDR_0_port );
   
   PC_REG : REG_GENERIC_NBIT32_0 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => PC_BUS_31_port, 
                           DATA_IN(30) => PC_BUS_30_port, DATA_IN(29) => 
                           PC_BUS_29_port, DATA_IN(28) => PC_BUS_28_port, 
                           DATA_IN(27) => PC_BUS_27_port, DATA_IN(26) => 
                           PC_BUS_26_port, DATA_IN(25) => PC_BUS_25_port, 
                           DATA_IN(24) => PC_BUS_24_port, DATA_IN(23) => 
                           PC_BUS_23_port, DATA_IN(22) => PC_BUS_22_port, 
                           DATA_IN(21) => PC_BUS_21_port, DATA_IN(20) => 
                           PC_BUS_20_port, DATA_IN(19) => PC_BUS_19_port, 
                           DATA_IN(18) => PC_BUS_18_port, DATA_IN(17) => 
                           PC_BUS_17_port, DATA_IN(16) => PC_BUS_16_port, 
                           DATA_IN(15) => PC_BUS_15_port, DATA_IN(14) => 
                           PC_BUS_14_port, DATA_IN(13) => PC_BUS_13_port, 
                           DATA_IN(12) => PC_BUS_12_port, DATA_IN(11) => 
                           PC_BUS_11_port, DATA_IN(10) => PC_BUS_10_port, 
                           DATA_IN(9) => PC_BUS_9_port, DATA_IN(8) => 
                           PC_BUS_8_port, DATA_IN(7) => PC_BUS_7_port, 
                           DATA_IN(6) => PC_BUS_6_port, DATA_IN(5) => 
                           PC_BUS_5_port, DATA_IN(4) => PC_BUS_4_port, 
                           DATA_IN(3) => PC_BUS_3_port, DATA_IN(2) => 
                           PC_BUS_2_port, DATA_IN(1) => PC_BUS_1_port, 
                           DATA_IN(0) => PC_BUS_0_port, DATA_OUT(31) => 
                           I_ADDR_31_port, DATA_OUT(30) => I_ADDR_30_port, 
                           DATA_OUT(29) => I_ADDR_29_port, DATA_OUT(28) => 
                           I_ADDR_28_port, DATA_OUT(27) => I_ADDR_27_port, 
                           DATA_OUT(26) => I_ADDR_26_port, DATA_OUT(25) => 
                           I_ADDR_25_port, DATA_OUT(24) => I_ADDR_24_port, 
                           DATA_OUT(23) => I_ADDR_23_port, DATA_OUT(22) => 
                           I_ADDR_22_port, DATA_OUT(21) => I_ADDR_21_port, 
                           DATA_OUT(20) => I_ADDR_20_port, DATA_OUT(19) => 
                           I_ADDR_19_port, DATA_OUT(18) => I_ADDR_18_port, 
                           DATA_OUT(17) => I_ADDR_17_port, DATA_OUT(16) => 
                           I_ADDR_16_port, DATA_OUT(15) => I_ADDR_15_port, 
                           DATA_OUT(14) => I_ADDR_14_port, DATA_OUT(13) => 
                           I_ADDR_13_port, DATA_OUT(12) => I_ADDR_12_port, 
                           DATA_OUT(11) => I_ADDR_11_port, DATA_OUT(10) => 
                           I_ADDR_10_port, DATA_OUT(9) => I_ADDR_9_port, 
                           DATA_OUT(8) => I_ADDR_8_port, DATA_OUT(7) => 
                           I_ADDR_7_port, DATA_OUT(6) => I_ADDR_6_port, 
                           DATA_OUT(5) => I_ADDR_5_port, DATA_OUT(4) => 
                           I_ADDR_4_port, DATA_OUT(3) => I_ADDR_3_port, 
                           DATA_OUT(2) => I_ADDR_2_port, DATA_OUT(1) => 
                           I_ADDR_1_port, DATA_OUT(0) => I_ADDR_0_port);
   DP : DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 port map( CLK => CLK
                           , RST => RST, IR_IN(31) => I_DATA(31), IR_IN(30) => 
                           I_DATA(30), IR_IN(29) => I_DATA(29), IR_IN(28) => 
                           I_DATA(28), IR_IN(27) => I_DATA(27), IR_IN(26) => 
                           I_DATA(26), IR_IN(25) => I_DATA(25), IR_IN(24) => 
                           I_DATA(24), IR_IN(23) => I_DATA(23), IR_IN(22) => 
                           I_DATA(22), IR_IN(21) => I_DATA(21), IR_IN(20) => 
                           I_DATA(20), IR_IN(19) => I_DATA(19), IR_IN(18) => 
                           I_DATA(18), IR_IN(17) => I_DATA(17), IR_IN(16) => 
                           I_DATA(16), IR_IN(15) => I_DATA(15), IR_IN(14) => 
                           I_DATA(14), IR_IN(13) => I_DATA(13), IR_IN(12) => 
                           I_DATA(12), IR_IN(11) => I_DATA(11), IR_IN(10) => 
                           I_DATA(10), IR_IN(9) => I_DATA(9), IR_IN(8) => 
                           I_DATA(8), IR_IN(7) => I_DATA(7), IR_IN(6) => 
                           I_DATA(6), IR_IN(5) => I_DATA(5), IR_IN(4) => 
                           I_DATA(4), IR_IN(3) => I_DATA(3), IR_IN(2) => 
                           I_DATA(2), IR_IN(1) => I_DATA(1), IR_IN(0) => 
                           I_DATA(0), IR_LATCH_EN => IR_LATCH_EN, NPC_LATCH_EN 
                           => NPC_LATCH_EN, RegA_LATCH_EN => RegA_LATCH_EN, 
                           RegB_LATCH_EN => RegB_LATCH_EN, RegIMM_LATCH_EN => 
                           RegIMM_LATCH_EN, SIGNED_IMM => SIGNED_IMM, MUXA_SEL 
                           => MUXA_SEL, MUXB_SEL => MUXB_SEL, ALU_OUTREG_EN => 
                           ALU_OUTREG_EN, EQ_COND => EQ_COND, IS_JUMP => 
                           IS_JUMP, ALU_OPCODE(0) => ALU_OPCODE_3_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_2_port, ALU_OPCODE(2) =>
                           ALU_OPCODE_1_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_0_port, JUMP_EN => JUMP_EN, PC_LATCH_EN 
                           => PC_LATCH_EN, IS_JAL => IS_JAL, WB_MUX_SEL => 
                           WB_MUX_SEL, RF_WE => RF_WE, D_ADDR(5) => D_ADDR(5), 
                           D_ADDR(4) => D_ADDR(4), D_ADDR(3) => D_ADDR(3), 
                           D_ADDR(2) => D_ADDR(2), D_ADDR(1) => D_ADDR(1), 
                           D_ADDR(0) => D_ADDR(0), D_DATA_IN(31) => 
                           D_DATA_IN(31), D_DATA_IN(30) => D_DATA_IN(30), 
                           D_DATA_IN(29) => D_DATA_IN(29), D_DATA_IN(28) => 
                           D_DATA_IN(28), D_DATA_IN(27) => D_DATA_IN(27), 
                           D_DATA_IN(26) => D_DATA_IN(26), D_DATA_IN(25) => 
                           D_DATA_IN(25), D_DATA_IN(24) => D_DATA_IN(24), 
                           D_DATA_IN(23) => D_DATA_IN(23), D_DATA_IN(22) => 
                           D_DATA_IN(22), D_DATA_IN(21) => D_DATA_IN(21), 
                           D_DATA_IN(20) => D_DATA_IN(20), D_DATA_IN(19) => 
                           D_DATA_IN(19), D_DATA_IN(18) => D_DATA_IN(18), 
                           D_DATA_IN(17) => D_DATA_IN(17), D_DATA_IN(16) => 
                           D_DATA_IN(16), D_DATA_IN(15) => D_DATA_IN(15), 
                           D_DATA_IN(14) => D_DATA_IN(14), D_DATA_IN(13) => 
                           D_DATA_IN(13), D_DATA_IN(12) => D_DATA_IN(12), 
                           D_DATA_IN(11) => D_DATA_IN(11), D_DATA_IN(10) => 
                           D_DATA_IN(10), D_DATA_IN(9) => D_DATA_IN(9), 
                           D_DATA_IN(8) => D_DATA_IN(8), D_DATA_IN(7) => 
                           D_DATA_IN(7), D_DATA_IN(6) => D_DATA_IN(6), 
                           D_DATA_IN(5) => D_DATA_IN(5), D_DATA_IN(4) => 
                           D_DATA_IN(4), D_DATA_IN(3) => D_DATA_IN(3), 
                           D_DATA_IN(2) => D_DATA_IN(2), D_DATA_IN(1) => 
                           D_DATA_IN(1), D_DATA_IN(0) => D_DATA_IN(0), 
                           D_DATA_OUT(31) => D_DATA_OUT(31), D_DATA_OUT(30) => 
                           D_DATA_OUT(30), D_DATA_OUT(29) => D_DATA_OUT(29), 
                           D_DATA_OUT(28) => D_DATA_OUT(28), D_DATA_OUT(27) => 
                           D_DATA_OUT(27), D_DATA_OUT(26) => D_DATA_OUT(26), 
                           D_DATA_OUT(25) => D_DATA_OUT(25), D_DATA_OUT(24) => 
                           D_DATA_OUT(24), D_DATA_OUT(23) => D_DATA_OUT(23), 
                           D_DATA_OUT(22) => D_DATA_OUT(22), D_DATA_OUT(21) => 
                           D_DATA_OUT(21), D_DATA_OUT(20) => D_DATA_OUT(20), 
                           D_DATA_OUT(19) => D_DATA_OUT(19), D_DATA_OUT(18) => 
                           D_DATA_OUT(18), D_DATA_OUT(17) => D_DATA_OUT(17), 
                           D_DATA_OUT(16) => D_DATA_OUT(16), D_DATA_OUT(15) => 
                           D_DATA_OUT(15), D_DATA_OUT(14) => D_DATA_OUT(14), 
                           D_DATA_OUT(13) => D_DATA_OUT(13), D_DATA_OUT(12) => 
                           D_DATA_OUT(12), D_DATA_OUT(11) => D_DATA_OUT(11), 
                           D_DATA_OUT(10) => D_DATA_OUT(10), D_DATA_OUT(9) => 
                           D_DATA_OUT(9), D_DATA_OUT(8) => D_DATA_OUT(8), 
                           D_DATA_OUT(7) => D_DATA_OUT(7), D_DATA_OUT(6) => 
                           D_DATA_OUT(6), D_DATA_OUT(5) => D_DATA_OUT(5), 
                           D_DATA_OUT(4) => D_DATA_OUT(4), D_DATA_OUT(3) => 
                           D_DATA_OUT(3), D_DATA_OUT(2) => D_DATA_OUT(2), 
                           D_DATA_OUT(1) => D_DATA_OUT(1), D_DATA_OUT(0) => 
                           D_DATA_OUT(0), PC_IN(31) => I_ADDR_31_port, 
                           PC_IN(30) => I_ADDR_30_port, PC_IN(29) => 
                           I_ADDR_29_port, PC_IN(28) => I_ADDR_28_port, 
                           PC_IN(27) => I_ADDR_27_port, PC_IN(26) => 
                           I_ADDR_26_port, PC_IN(25) => I_ADDR_25_port, 
                           PC_IN(24) => I_ADDR_24_port, PC_IN(23) => 
                           I_ADDR_23_port, PC_IN(22) => I_ADDR_22_port, 
                           PC_IN(21) => I_ADDR_21_port, PC_IN(20) => 
                           I_ADDR_20_port, PC_IN(19) => I_ADDR_19_port, 
                           PC_IN(18) => I_ADDR_18_port, PC_IN(17) => 
                           I_ADDR_17_port, PC_IN(16) => I_ADDR_16_port, 
                           PC_IN(15) => I_ADDR_15_port, PC_IN(14) => 
                           I_ADDR_14_port, PC_IN(13) => I_ADDR_13_port, 
                           PC_IN(12) => I_ADDR_12_port, PC_IN(11) => 
                           I_ADDR_11_port, PC_IN(10) => I_ADDR_10_port, 
                           PC_IN(9) => I_ADDR_9_port, PC_IN(8) => I_ADDR_8_port
                           , PC_IN(7) => I_ADDR_7_port, PC_IN(6) => 
                           I_ADDR_6_port, PC_IN(5) => I_ADDR_5_port, PC_IN(4) 
                           => I_ADDR_4_port, PC_IN(3) => I_ADDR_3_port, 
                           PC_IN(2) => I_ADDR_2_port, PC_IN(1) => I_ADDR_1_port
                           , PC_IN(0) => I_ADDR_0_port, PC_BUS(31) => 
                           PC_BUS_31_port, PC_BUS(30) => PC_BUS_30_port, 
                           PC_BUS(29) => PC_BUS_29_port, PC_BUS(28) => 
                           PC_BUS_28_port, PC_BUS(27) => PC_BUS_27_port, 
                           PC_BUS(26) => PC_BUS_26_port, PC_BUS(25) => 
                           PC_BUS_25_port, PC_BUS(24) => PC_BUS_24_port, 
                           PC_BUS(23) => PC_BUS_23_port, PC_BUS(22) => 
                           PC_BUS_22_port, PC_BUS(21) => PC_BUS_21_port, 
                           PC_BUS(20) => PC_BUS_20_port, PC_BUS(19) => 
                           PC_BUS_19_port, PC_BUS(18) => PC_BUS_18_port, 
                           PC_BUS(17) => PC_BUS_17_port, PC_BUS(16) => 
                           PC_BUS_16_port, PC_BUS(15) => PC_BUS_15_port, 
                           PC_BUS(14) => PC_BUS_14_port, PC_BUS(13) => 
                           PC_BUS_13_port, PC_BUS(12) => PC_BUS_12_port, 
                           PC_BUS(11) => PC_BUS_11_port, PC_BUS(10) => 
                           PC_BUS_10_port, PC_BUS(9) => PC_BUS_9_port, 
                           PC_BUS(8) => PC_BUS_8_port, PC_BUS(7) => 
                           PC_BUS_7_port, PC_BUS(6) => PC_BUS_6_port, PC_BUS(5)
                           => PC_BUS_5_port, PC_BUS(4) => PC_BUS_4_port, 
                           PC_BUS(3) => PC_BUS_3_port, PC_BUS(2) => 
                           PC_BUS_2_port, PC_BUS(1) => PC_BUS_1_port, PC_BUS(0)
                           => PC_BUS_0_port);
   CU : dlx_cu port map( Clk => CLK, Rst => RST, IR_IN(31) => I_DATA(31), 
                           IR_IN(30) => I_DATA(30), IR_IN(29) => I_DATA(29), 
                           IR_IN(28) => I_DATA(28), IR_IN(27) => I_DATA(27), 
                           IR_IN(26) => I_DATA(26), IR_IN(25) => I_DATA(25), 
                           IR_IN(24) => I_DATA(24), IR_IN(23) => I_DATA(23), 
                           IR_IN(22) => I_DATA(22), IR_IN(21) => I_DATA(21), 
                           IR_IN(20) => I_DATA(20), IR_IN(19) => I_DATA(19), 
                           IR_IN(18) => I_DATA(18), IR_IN(17) => I_DATA(17), 
                           IR_IN(16) => I_DATA(16), IR_IN(15) => I_DATA(15), 
                           IR_IN(14) => I_DATA(14), IR_IN(13) => I_DATA(13), 
                           IR_IN(12) => I_DATA(12), IR_IN(11) => I_DATA(11), 
                           IR_IN(10) => I_DATA(10), IR_IN(9) => I_DATA(9), 
                           IR_IN(8) => I_DATA(8), IR_IN(7) => I_DATA(7), 
                           IR_IN(6) => I_DATA(6), IR_IN(5) => I_DATA(5), 
                           IR_IN(4) => I_DATA(4), IR_IN(3) => I_DATA(3), 
                           IR_IN(2) => I_DATA(2), IR_IN(1) => I_DATA(1), 
                           IR_IN(0) => I_DATA(0), IR_LATCH_EN => n_2158, 
                           NPC_LATCH_EN => n_2159, RegA_LATCH_EN => n_2160, 
                           RegB_LATCH_EN => n_2161, RegIMM_LATCH_EN => n_2162, 
                           SIGNED_IMM => n_2163, MUXA_SEL => n_2164, MUXB_SEL 
                           => n_2165, ALU_OUTREG_EN => n_2166, EQ_COND => 
                           n_2167, IS_JUMP => n_2168, ALU_OPCODE(0) => 
                           ALU_OPCODE_3_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_2_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_1_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_0_port, DRAM_WE => n_2169, LMD_LATCH_EN 
                           => n_2170, JUMP_EN => n_2171, PC_LATCH_EN => n_2172,
                           IS_JAL => n_2173, WB_MUX_SEL => n_2174, RF_WE => 
                           n_2175);
   RF_WE <= '0';
   WB_MUX_SEL <= '0';
   IS_JAL <= '0';
   PC_LATCH_EN <= '0';
   JUMP_EN <= '0';
   D_RR <= '0';
   D_WR <= '0';
   IS_JUMP <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   SIGNED_IMM <= '0';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   NPC_LATCH_EN <= '0';
   IR_LATCH_EN <= '0';

end SYN_DLX_RTL;

library IEEE;

use IEEE.std_logic_1164.all;
entity SELECT_OP is
   generic ( num_inputs, input_width : integer );
   port(
      DATA : in std_logic_vector( num_inputs  * input_width - 1 downto 0 );
      CONTROL : in std_logic_vector( num_inputs - 1 downto 0 );
      Z : out std_logic_vector( input_width - 1 downto 0 )
   );
end SELECT_OP;

architecture RTL of SELECT_OP is
begin

   process ( DATA, CONTROL )
      variable index, high, low : integer;
   begin
   
      --  Initialize variables
      index := 0;
      
      -- Loop over the values of the control inputs
      for_loop : for i in CONTROL'range loop
      
         if ( CONTROL(i) = '1' ) then
         
            index := i;
            exit for_loop;
            
         end if;
         
      end loop;
      
      -- Store the corresponding data lines into the output
      low := input_width * index;
      high := low + input_width - 1;
      Z <= DATA( high downto low );
   
   end process;
   
end RTL;

library IEEE;

use IEEE.std_logic_1164.all;

entity SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT is
   generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
   port(
      clear, preset, enable, data_in, synch_clear, synch_preset, synch_toggle, 
         synch_enable, next_state, clocked_on : in std_logic;
      Q, QN : buffer std_logic
   );
end SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT;

architecture RTL of SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT is
begin

   process ( preset, clear, enable, data_in, clocked_on )
   begin
   
            -- Check the value of inputs (asynchronous first)
            if ( ( ( preset /= '1' ) and ( preset /= '0' ) ) or ( ( clear /= 
                     '1' ) and ( clear /= '0' ) )  ) then
               Q <= 'X';
            elsif ( clear = '1' and preset = '1' ) then
               case ac_as_q is
                  when 2 =>
                     Q <= '1';
                  when 1 =>
                     Q <= '0';
                  when others =>
                     Q <= 'X';
               end case;
               case ac_as_qn is
                  when 2 =>
                     QN <= '1';
                  when 1 =>
                     QN <= '0';
                  when others =>
                     QN <= 'X';
               end case;
            elsif ( clear = '1' ) then
               Q <= '0';
            elsif ( preset = '1' ) then
               Q <= '1';
            elsif ( ( enable /= '1' ) and ( enable /= '0' ) ) then
               Q <= 'X';
            elsif ( enable = '1' ) then
               Q <= data_in;
            elsif ( ( clocked_on /= '1' ) and ( clocked_on /= '0' ) ) then
               Q <= 'X';
            elsif ( clocked_on'event and clocked_on = '1' ) then
         if ( ( ( synch_preset /= '1' ) and ( synch_preset /= '0' ) ) or ( ( 
                  synch_clear /= '1' ) and ( synch_clear /= '0' ) )  ) then
            Q <= 'X';
         elsif ( synch_clear = '1' and synch_preset = '1' ) then
            case sc_ss_q is
               when 2 =>
                  Q <= '1';
               when 1 =>
                  Q <= '0';
               when others =>
                  Q <= 'X';
            end case;
         elsif ( synch_clear = '1' ) then
            Q <= '0';
         elsif ( synch_preset = '1' ) then
            Q <= '1';
         elsif ( ( ( synch_toggle /= '1' ) and ( synch_toggle /= '0' ) ) or ( (
                  synch_enable /= '1' ) and ( synch_enable /= '0' ) )  ) then
            Q <= 'X';
         elsif ( synch_enable = '1' and synch_toggle = '1' ) then
            Q <= 'X';
         elsif ( synch_toggle = '1' ) then
            Q <= QN;
         elsif ( synch_enable = '1' ) then
            Q <= next_state;
         end if;
      end if;
   
   end process;

end RTL;
