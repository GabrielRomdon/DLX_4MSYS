
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOpType is (NOP, ADDS, SUBS, ANDS, ORS, XORS, SLE, SGE, SNE, SRLS, SLLS)
   ;
attribute ENUM_ENCODING of aluOpType : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOpType(arg : in std_logic_vector( 1 to 4 )) 
               return aluOpType;
   function aluOpType_to_std_logic_vector(arg : in aluOpType) return 
               std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOpType(arg : in std_logic_vector( 1 to 4 )) 
   return aluOpType is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "0000" => return NOP;
         when "0001" => return ADDS;
         when "0010" => return SUBS;
         when "0011" => return ANDS;
         when "0100" => return ORS;
         when "0101" => return XORS;
         when "0110" => return SLE;
         when "0111" => return SGE;
         when "1000" => return SNE;
         when "1001" => return SRLS;
         when "1010" => return SLLS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOpType_to_std_logic_vector(arg : in aluOpType) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "0000";
         when ADDS => return "0001";
         when SUBS => return "0010";
         when ANDS => return "0011";
         when ORS => return "0100";
         when XORS => return "0101";
         when SLE => return "0110";
         when SGE => return "0111";
         when SNE => return "1000";
         when SRLS => return "1001";
         when SLLS => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_127 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_127;

architecture SYN_BEHAVIOUR of NAND3_127 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_126 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_126;

architecture SYN_BEHAVIOUR of NAND3_126 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_125 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_125;

architecture SYN_BEHAVIOUR of NAND3_125 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_124 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_124;

architecture SYN_BEHAVIOUR of NAND3_124 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_123 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_123;

architecture SYN_BEHAVIOUR of NAND3_123 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_122 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_122;

architecture SYN_BEHAVIOUR of NAND3_122 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_121 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_121;

architecture SYN_BEHAVIOUR of NAND3_121 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_120 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_120;

architecture SYN_BEHAVIOUR of NAND3_120 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_119 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_119;

architecture SYN_BEHAVIOUR of NAND3_119 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_118 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_118;

architecture SYN_BEHAVIOUR of NAND3_118 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_117 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_117;

architecture SYN_BEHAVIOUR of NAND3_117 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_116 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_116;

architecture SYN_BEHAVIOUR of NAND3_116 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_115 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_115;

architecture SYN_BEHAVIOUR of NAND3_115 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_114 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_114;

architecture SYN_BEHAVIOUR of NAND3_114 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_113 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_113;

architecture SYN_BEHAVIOUR of NAND3_113 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_112 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_112;

architecture SYN_BEHAVIOUR of NAND3_112 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_111 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_111;

architecture SYN_BEHAVIOUR of NAND3_111 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_110 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_110;

architecture SYN_BEHAVIOUR of NAND3_110 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_109 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_109;

architecture SYN_BEHAVIOUR of NAND3_109 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_108 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_108;

architecture SYN_BEHAVIOUR of NAND3_108 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_107 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_107;

architecture SYN_BEHAVIOUR of NAND3_107 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_106 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_106;

architecture SYN_BEHAVIOUR of NAND3_106 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_105 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_105;

architecture SYN_BEHAVIOUR of NAND3_105 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_104 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_104;

architecture SYN_BEHAVIOUR of NAND3_104 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_103 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_103;

architecture SYN_BEHAVIOUR of NAND3_103 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_102 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_102;

architecture SYN_BEHAVIOUR of NAND3_102 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_101 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_101;

architecture SYN_BEHAVIOUR of NAND3_101 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_100 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_100;

architecture SYN_BEHAVIOUR of NAND3_100 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_99 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_99;

architecture SYN_BEHAVIOUR of NAND3_99 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_98 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_98;

architecture SYN_BEHAVIOUR of NAND3_98 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_97 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_97;

architecture SYN_BEHAVIOUR of NAND3_97 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_31 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_31;

architecture SYN_BEHAVIOUR of NAND4_31 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_30 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_30;

architecture SYN_BEHAVIOUR of NAND4_30 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_29 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_29;

architecture SYN_BEHAVIOUR of NAND4_29 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_28 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_28;

architecture SYN_BEHAVIOUR of NAND4_28 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_27 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_27;

architecture SYN_BEHAVIOUR of NAND4_27 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_26 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_26;

architecture SYN_BEHAVIOUR of NAND4_26 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_25 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_25;

architecture SYN_BEHAVIOUR of NAND4_25 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_24 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_24;

architecture SYN_BEHAVIOUR of NAND4_24 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_23 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_23;

architecture SYN_BEHAVIOUR of NAND4_23 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_22 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_22;

architecture SYN_BEHAVIOUR of NAND4_22 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_21 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_21;

architecture SYN_BEHAVIOUR of NAND4_21 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_20 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_20;

architecture SYN_BEHAVIOUR of NAND4_20 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_19 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_19;

architecture SYN_BEHAVIOUR of NAND4_19 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_18 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_18;

architecture SYN_BEHAVIOUR of NAND4_18 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_17 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_17;

architecture SYN_BEHAVIOUR of NAND4_17 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_16 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_16;

architecture SYN_BEHAVIOUR of NAND4_16 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_15 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_15;

architecture SYN_BEHAVIOUR of NAND4_15 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_14 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_14;

architecture SYN_BEHAVIOUR of NAND4_14 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_13 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_13;

architecture SYN_BEHAVIOUR of NAND4_13 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_12 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_12;

architecture SYN_BEHAVIOUR of NAND4_12 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_11 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_11;

architecture SYN_BEHAVIOUR of NAND4_11 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_10 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_10;

architecture SYN_BEHAVIOUR of NAND4_10 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_9 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_9;

architecture SYN_BEHAVIOUR of NAND4_9 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_8 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_8;

architecture SYN_BEHAVIOUR of NAND4_8 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_7 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_7;

architecture SYN_BEHAVIOUR of NAND4_7 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_6 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_6;

architecture SYN_BEHAVIOUR of NAND4_6 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_5 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_5;

architecture SYN_BEHAVIOUR of NAND4_5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_4 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_4;

architecture SYN_BEHAVIOUR of NAND4_4 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_3 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_3;

architecture SYN_BEHAVIOUR of NAND4_3 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_2 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_2;

architecture SYN_BEHAVIOUR of NAND4_2 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_1 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_1;

architecture SYN_BEHAVIOUR of NAND4_1 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_95 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_95;

architecture SYN_BEHAVIOUR of NAND3_95 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_94 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_94;

architecture SYN_BEHAVIOUR of NAND3_94 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_93 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_93;

architecture SYN_BEHAVIOUR of NAND3_93 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_92 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_92;

architecture SYN_BEHAVIOUR of NAND3_92 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_91 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_91;

architecture SYN_BEHAVIOUR of NAND3_91 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_90 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_90;

architecture SYN_BEHAVIOUR of NAND3_90 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_89 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_89;

architecture SYN_BEHAVIOUR of NAND3_89 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_88 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_88;

architecture SYN_BEHAVIOUR of NAND3_88 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_87 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_87;

architecture SYN_BEHAVIOUR of NAND3_87 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_86 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_86;

architecture SYN_BEHAVIOUR of NAND3_86 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_85 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_85;

architecture SYN_BEHAVIOUR of NAND3_85 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_84 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_84;

architecture SYN_BEHAVIOUR of NAND3_84 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_83 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_83;

architecture SYN_BEHAVIOUR of NAND3_83 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_82 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_82;

architecture SYN_BEHAVIOUR of NAND3_82 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_81 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_81;

architecture SYN_BEHAVIOUR of NAND3_81 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_80 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_80;

architecture SYN_BEHAVIOUR of NAND3_80 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_79 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_79;

architecture SYN_BEHAVIOUR of NAND3_79 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_78 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_78;

architecture SYN_BEHAVIOUR of NAND3_78 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_77 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_77;

architecture SYN_BEHAVIOUR of NAND3_77 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_76 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_76;

architecture SYN_BEHAVIOUR of NAND3_76 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_75 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_75;

architecture SYN_BEHAVIOUR of NAND3_75 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_74 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_74;

architecture SYN_BEHAVIOUR of NAND3_74 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_73 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_73;

architecture SYN_BEHAVIOUR of NAND3_73 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_72 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_72;

architecture SYN_BEHAVIOUR of NAND3_72 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_71 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_71;

architecture SYN_BEHAVIOUR of NAND3_71 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_70 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_70;

architecture SYN_BEHAVIOUR of NAND3_70 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_69 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_69;

architecture SYN_BEHAVIOUR of NAND3_69 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_68 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_68;

architecture SYN_BEHAVIOUR of NAND3_68 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_67 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_67;

architecture SYN_BEHAVIOUR of NAND3_67 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_66 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_66;

architecture SYN_BEHAVIOUR of NAND3_66 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_65 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_65;

architecture SYN_BEHAVIOUR of NAND3_65 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_64 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_64;

architecture SYN_BEHAVIOUR of NAND3_64 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_63 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_63;

architecture SYN_BEHAVIOUR of NAND3_63 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_62 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_62;

architecture SYN_BEHAVIOUR of NAND3_62 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_61 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_61;

architecture SYN_BEHAVIOUR of NAND3_61 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_60 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_60;

architecture SYN_BEHAVIOUR of NAND3_60 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_59 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_59;

architecture SYN_BEHAVIOUR of NAND3_59 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_58 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_58;

architecture SYN_BEHAVIOUR of NAND3_58 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_57 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_57;

architecture SYN_BEHAVIOUR of NAND3_57 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_56 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_56;

architecture SYN_BEHAVIOUR of NAND3_56 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_55 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_55;

architecture SYN_BEHAVIOUR of NAND3_55 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_54 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_54;

architecture SYN_BEHAVIOUR of NAND3_54 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_53 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_53;

architecture SYN_BEHAVIOUR of NAND3_53 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_52 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_52;

architecture SYN_BEHAVIOUR of NAND3_52 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_51 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_51;

architecture SYN_BEHAVIOUR of NAND3_51 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_50 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_50;

architecture SYN_BEHAVIOUR of NAND3_50 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_49 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_49;

architecture SYN_BEHAVIOUR of NAND3_49 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_48 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_48;

architecture SYN_BEHAVIOUR of NAND3_48 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_47 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_47;

architecture SYN_BEHAVIOUR of NAND3_47 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_46 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_46;

architecture SYN_BEHAVIOUR of NAND3_46 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_45 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_45;

architecture SYN_BEHAVIOUR of NAND3_45 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_44 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_44;

architecture SYN_BEHAVIOUR of NAND3_44 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_43 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_43;

architecture SYN_BEHAVIOUR of NAND3_43 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_42 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_42;

architecture SYN_BEHAVIOUR of NAND3_42 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_41 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_41;

architecture SYN_BEHAVIOUR of NAND3_41 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_40 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_40;

architecture SYN_BEHAVIOUR of NAND3_40 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_39 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_39;

architecture SYN_BEHAVIOUR of NAND3_39 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_38 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_38;

architecture SYN_BEHAVIOUR of NAND3_38 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_37 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_37;

architecture SYN_BEHAVIOUR of NAND3_37 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_36 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_36;

architecture SYN_BEHAVIOUR of NAND3_36 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_35 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_35;

architecture SYN_BEHAVIOUR of NAND3_35 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_34 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_34;

architecture SYN_BEHAVIOUR of NAND3_34 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_33 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_33;

architecture SYN_BEHAVIOUR of NAND3_33 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_32 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_32;

architecture SYN_BEHAVIOUR of NAND3_32 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_31 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_31;

architecture SYN_BEHAVIOUR of NAND3_31 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_30 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_30;

architecture SYN_BEHAVIOUR of NAND3_30 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_29 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_29;

architecture SYN_BEHAVIOUR of NAND3_29 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_28 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_28;

architecture SYN_BEHAVIOUR of NAND3_28 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_27 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_27;

architecture SYN_BEHAVIOUR of NAND3_27 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_26 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_26;

architecture SYN_BEHAVIOUR of NAND3_26 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_25 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_25;

architecture SYN_BEHAVIOUR of NAND3_25 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_24 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_24;

architecture SYN_BEHAVIOUR of NAND3_24 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_23 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_23;

architecture SYN_BEHAVIOUR of NAND3_23 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_22 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_22;

architecture SYN_BEHAVIOUR of NAND3_22 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_21 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_21;

architecture SYN_BEHAVIOUR of NAND3_21 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_20 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_20;

architecture SYN_BEHAVIOUR of NAND3_20 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_19 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_19;

architecture SYN_BEHAVIOUR of NAND3_19 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_18 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_18;

architecture SYN_BEHAVIOUR of NAND3_18 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_17 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_17;

architecture SYN_BEHAVIOUR of NAND3_17 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_16 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_16;

architecture SYN_BEHAVIOUR of NAND3_16 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_15 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_15;

architecture SYN_BEHAVIOUR of NAND3_15 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_14 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_14;

architecture SYN_BEHAVIOUR of NAND3_14 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_13 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_13;

architecture SYN_BEHAVIOUR of NAND3_13 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_12 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_12;

architecture SYN_BEHAVIOUR of NAND3_12 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_11 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_11;

architecture SYN_BEHAVIOUR of NAND3_11 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_10 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_10;

architecture SYN_BEHAVIOUR of NAND3_10 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_9 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_9;

architecture SYN_BEHAVIOUR of NAND3_9 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_8 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_8;

architecture SYN_BEHAVIOUR of NAND3_8 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_7 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_7;

architecture SYN_BEHAVIOUR of NAND3_7 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_6 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_6;

architecture SYN_BEHAVIOUR of NAND3_6 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_5 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_5;

architecture SYN_BEHAVIOUR of NAND3_5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_4 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_4;

architecture SYN_BEHAVIOUR of NAND3_4 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_3 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_3;

architecture SYN_BEHAVIOUR of NAND3_3 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_2 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_2;

architecture SYN_BEHAVIOUR of NAND3_2 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_1 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_1;

architecture SYN_BEHAVIOUR of NAND3_1 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_1;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT5_1 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 downto 
         0);  DATA_OUT : out std_logic_vector (4 downto 0));

end REG_GENERIC_NBIT5_1;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n9, n14, n15, n16, n17, n18, n19
      , n_1000, n_1001, n_1002, n_1003, n_1004 : std_logic;

begin
   DATA_OUT <= ( DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, 
      DATA_OUT_1_port, DATA_OUT_0_port );
   
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n3, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_1000);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n4, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_1001);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n5, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_1002);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n6, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_1003);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n9, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_1004);
   U7 : AOI22_X1 port map( A1 => DATA_IN(4), A2 => n18, B1 => DATA_OUT_4_port, 
                           B2 => n1, ZN => n14);
   U6 : AOI22_X1 port map( A1 => DATA_IN(3), A2 => n18, B1 => DATA_OUT_3_port, 
                           B2 => n1, ZN => n15);
   U5 : AOI22_X1 port map( A1 => DATA_IN(2), A2 => n18, B1 => DATA_OUT_2_port, 
                           B2 => n1, ZN => n16);
   U4 : AOI22_X1 port map( A1 => DATA_IN(1), A2 => n18, B1 => DATA_OUT_1_port, 
                           B2 => n1, ZN => n17);
   U3 : AOI22_X1 port map( A1 => DATA_IN(0), A2 => n18, B1 => DATA_OUT_0_port, 
                           B2 => n1, ZN => n19);
   U8 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => n18);
   U9 : NOR2_X1 port map( A1 => EN, A2 => n2, ZN => n1);
   U10 : INV_X1 port map( A => RST, ZN => n2);
   U11 : INV_X1 port map( A => n19, ZN => n9);
   U12 : INV_X1 port map( A => n17, ZN => n6);
   U13 : INV_X1 port map( A => n16, ZN => n5);
   U14 : INV_X1 port map( A => n15, ZN => n4);
   U15 : INV_X1 port map( A => n14, ZN => n3);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_7 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_7;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036 : 
      std_logic;

begin
   DATA_OUT <= ( DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port );
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n44, CK => CLK, Q => 
                           DATA_OUT_31_port, QN => n_1005);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n45, CK => CLK, Q => 
                           DATA_OUT_30_port, QN => n_1006);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n46, CK => CLK, Q => 
                           DATA_OUT_29_port, QN => n_1007);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n47, CK => CLK, Q => 
                           DATA_OUT_28_port, QN => n_1008);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n48, CK => CLK, Q => 
                           DATA_OUT_27_port, QN => n_1009);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n49, CK => CLK, Q => 
                           DATA_OUT_26_port, QN => n_1010);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n50, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_1011);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n51, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n_1012);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n52, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_1013);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n53, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n_1014);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n54, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n_1015);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n55, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_1016);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n56, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_1017);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n57, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_1018);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n58, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_1019);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n59, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n_1020);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n60, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n_1021);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n61, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n_1022);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n62, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n_1023);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n63, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n_1024);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n64, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n_1025);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n65, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n_1026);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n66, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n_1027);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n67, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n_1028);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n_1029);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n_1030);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT_5_port, QN => n_1031);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_1032);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_1033);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_1034);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_1035);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_1036);
   U3 : BUF_X2 port map( A => n42, Z => n7);
   U4 : BUF_X2 port map( A => n42, Z => n8);
   U5 : BUF_X1 port map( A => n1, Z => n4);
   U6 : BUF_X1 port map( A => n1, Z => n5);
   U7 : BUF_X1 port map( A => n42, Z => n9);
   U8 : BUF_X1 port map( A => n1, Z => n6);
   U9 : AND2_X1 port map( A1 => n2, A2 => n10, ZN => n1);
   U10 : INV_X1 port map( A => n3, ZN => n2);
   U11 : INV_X1 port map( A => RST, ZN => n3);
   U12 : OR2_X1 port map( A1 => EN, A2 => n3, ZN => n10);
   U13 : INV_X1 port map( A => n10, ZN => n42);
   U14 : AOI22_X1 port map( A1 => DATA_OUT_0_port, A2 => n7, B1 => DATA_IN(0), 
                           B2 => n4, ZN => n11);
   U15 : INV_X1 port map( A => n11, ZN => n75);
   U16 : AOI22_X1 port map( A1 => DATA_OUT_1_port, A2 => n7, B1 => DATA_IN(1), 
                           B2 => n4, ZN => n12);
   U17 : INV_X1 port map( A => n12, ZN => n74);
   U18 : AOI22_X1 port map( A1 => DATA_OUT_2_port, A2 => n7, B1 => DATA_IN(2), 
                           B2 => n4, ZN => n13);
   U19 : INV_X1 port map( A => n13, ZN => n73);
   U20 : AOI22_X1 port map( A1 => DATA_OUT_3_port, A2 => n7, B1 => DATA_IN(3), 
                           B2 => n4, ZN => n14);
   U21 : INV_X1 port map( A => n14, ZN => n72);
   U22 : AOI22_X1 port map( A1 => DATA_OUT_4_port, A2 => n7, B1 => DATA_IN(4), 
                           B2 => n4, ZN => n15);
   U23 : INV_X1 port map( A => n15, ZN => n71);
   U24 : AOI22_X1 port map( A1 => DATA_OUT_5_port, A2 => n7, B1 => DATA_IN(5), 
                           B2 => n4, ZN => n16);
   U25 : INV_X1 port map( A => n16, ZN => n70);
   U26 : AOI22_X1 port map( A1 => DATA_OUT_6_port, A2 => n7, B1 => DATA_IN(6), 
                           B2 => n4, ZN => n17);
   U27 : INV_X1 port map( A => n17, ZN => n69);
   U28 : AOI22_X1 port map( A1 => DATA_OUT_7_port, A2 => n7, B1 => DATA_IN(7), 
                           B2 => n4, ZN => n18);
   U29 : INV_X1 port map( A => n18, ZN => n68);
   U30 : AOI22_X1 port map( A1 => DATA_OUT_8_port, A2 => n7, B1 => DATA_IN(8), 
                           B2 => n4, ZN => n19);
   U31 : INV_X1 port map( A => n19, ZN => n67);
   U32 : AOI22_X1 port map( A1 => DATA_OUT_9_port, A2 => n7, B1 => DATA_IN(9), 
                           B2 => n4, ZN => n20);
   U33 : INV_X1 port map( A => n20, ZN => n66);
   U34 : AOI22_X1 port map( A1 => DATA_OUT_10_port, A2 => n7, B1 => DATA_IN(10)
                           , B2 => n4, ZN => n21);
   U35 : INV_X1 port map( A => n21, ZN => n65);
   U36 : AOI22_X1 port map( A1 => DATA_OUT_11_port, A2 => n7, B1 => DATA_IN(11)
                           , B2 => n4, ZN => n22);
   U37 : INV_X1 port map( A => n22, ZN => n64);
   U38 : AOI22_X1 port map( A1 => DATA_OUT_12_port, A2 => n8, B1 => DATA_IN(12)
                           , B2 => n5, ZN => n23);
   U39 : INV_X1 port map( A => n23, ZN => n63);
   U40 : AOI22_X1 port map( A1 => DATA_OUT_13_port, A2 => n8, B1 => DATA_IN(13)
                           , B2 => n5, ZN => n24);
   U41 : INV_X1 port map( A => n24, ZN => n62);
   U42 : AOI22_X1 port map( A1 => DATA_OUT_14_port, A2 => n8, B1 => DATA_IN(14)
                           , B2 => n5, ZN => n25);
   U43 : INV_X1 port map( A => n25, ZN => n61);
   U44 : AOI22_X1 port map( A1 => DATA_OUT_15_port, A2 => n8, B1 => DATA_IN(15)
                           , B2 => n5, ZN => n26);
   U45 : INV_X1 port map( A => n26, ZN => n60);
   U46 : AOI22_X1 port map( A1 => DATA_OUT_16_port, A2 => n8, B1 => DATA_IN(16)
                           , B2 => n5, ZN => n27);
   U47 : INV_X1 port map( A => n27, ZN => n59);
   U48 : AOI22_X1 port map( A1 => DATA_OUT_17_port, A2 => n8, B1 => DATA_IN(17)
                           , B2 => n5, ZN => n28);
   U49 : INV_X1 port map( A => n28, ZN => n58);
   U50 : AOI22_X1 port map( A1 => DATA_OUT_18_port, A2 => n8, B1 => DATA_IN(18)
                           , B2 => n5, ZN => n29);
   U51 : INV_X1 port map( A => n29, ZN => n57);
   U52 : AOI22_X1 port map( A1 => DATA_OUT_19_port, A2 => n8, B1 => DATA_IN(19)
                           , B2 => n5, ZN => n30);
   U53 : INV_X1 port map( A => n30, ZN => n56);
   U54 : AOI22_X1 port map( A1 => DATA_OUT_20_port, A2 => n8, B1 => DATA_IN(20)
                           , B2 => n5, ZN => n31);
   U55 : INV_X1 port map( A => n31, ZN => n55);
   U56 : AOI22_X1 port map( A1 => DATA_OUT_21_port, A2 => n8, B1 => DATA_IN(21)
                           , B2 => n5, ZN => n32);
   U57 : INV_X1 port map( A => n32, ZN => n54);
   U58 : AOI22_X1 port map( A1 => DATA_OUT_22_port, A2 => n8, B1 => DATA_IN(22)
                           , B2 => n5, ZN => n33);
   U59 : INV_X1 port map( A => n33, ZN => n53);
   U60 : AOI22_X1 port map( A1 => DATA_OUT_23_port, A2 => n8, B1 => DATA_IN(23)
                           , B2 => n5, ZN => n34);
   U61 : INV_X1 port map( A => n34, ZN => n52);
   U62 : AOI22_X1 port map( A1 => DATA_OUT_24_port, A2 => n9, B1 => DATA_IN(24)
                           , B2 => n6, ZN => n35);
   U63 : INV_X1 port map( A => n35, ZN => n51);
   U64 : AOI22_X1 port map( A1 => DATA_OUT_25_port, A2 => n9, B1 => DATA_IN(25)
                           , B2 => n6, ZN => n36);
   U65 : INV_X1 port map( A => n36, ZN => n50);
   U66 : AOI22_X1 port map( A1 => DATA_OUT_26_port, A2 => n9, B1 => DATA_IN(26)
                           , B2 => n6, ZN => n37);
   U67 : INV_X1 port map( A => n37, ZN => n49);
   U68 : AOI22_X1 port map( A1 => DATA_OUT_27_port, A2 => n9, B1 => DATA_IN(27)
                           , B2 => n6, ZN => n38);
   U69 : INV_X1 port map( A => n38, ZN => n48);
   U70 : AOI22_X1 port map( A1 => DATA_OUT_28_port, A2 => n9, B1 => DATA_IN(28)
                           , B2 => n6, ZN => n39);
   U71 : INV_X1 port map( A => n39, ZN => n47);
   U72 : AOI22_X1 port map( A1 => DATA_OUT_29_port, A2 => n9, B1 => DATA_IN(29)
                           , B2 => n6, ZN => n40);
   U73 : INV_X1 port map( A => n40, ZN => n46);
   U74 : AOI22_X1 port map( A1 => DATA_OUT_30_port, A2 => n9, B1 => DATA_IN(30)
                           , B2 => n6, ZN => n41);
   U75 : INV_X1 port map( A => n41, ZN => n45);
   U76 : AOI22_X1 port map( A1 => DATA_OUT_31_port, A2 => n9, B1 => DATA_IN(31)
                           , B2 => n6, ZN => n43);
   U77 : INV_X1 port map( A => n43, ZN => n44);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_6 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_6;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068 : 
      std_logic;

begin
   DATA_OUT <= ( DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port );
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n44, CK => CLK, Q => 
                           DATA_OUT_31_port, QN => n_1037);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n45, CK => CLK, Q => 
                           DATA_OUT_30_port, QN => n_1038);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n46, CK => CLK, Q => 
                           DATA_OUT_29_port, QN => n_1039);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n47, CK => CLK, Q => 
                           DATA_OUT_28_port, QN => n_1040);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n48, CK => CLK, Q => 
                           DATA_OUT_27_port, QN => n_1041);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n49, CK => CLK, Q => 
                           DATA_OUT_26_port, QN => n_1042);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n50, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_1043);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n51, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n_1044);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n52, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_1045);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n53, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n_1046);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n54, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n_1047);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n55, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_1048);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n56, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_1049);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n57, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_1050);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n58, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_1051);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n59, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n_1052);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n60, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n_1053);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n61, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n_1054);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n62, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n_1055);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n63, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n_1056);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n64, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n_1057);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n65, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n_1058);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n66, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n_1059);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n67, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n_1060);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n_1061);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n_1062);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT_5_port, QN => n_1063);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_1064);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_1065);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_1066);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_1067);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_1068);
   U3 : BUF_X2 port map( A => n42, Z => n7);
   U4 : BUF_X2 port map( A => n42, Z => n8);
   U5 : BUF_X1 port map( A => n1, Z => n4);
   U6 : BUF_X1 port map( A => n1, Z => n5);
   U7 : BUF_X1 port map( A => n42, Z => n9);
   U8 : BUF_X1 port map( A => n1, Z => n6);
   U9 : AND2_X1 port map( A1 => n2, A2 => n10, ZN => n1);
   U10 : INV_X1 port map( A => n3, ZN => n2);
   U11 : INV_X1 port map( A => RST, ZN => n3);
   U12 : OR2_X1 port map( A1 => EN, A2 => n3, ZN => n10);
   U13 : INV_X1 port map( A => n10, ZN => n42);
   U14 : AOI22_X1 port map( A1 => DATA_OUT_0_port, A2 => n7, B1 => DATA_IN(0), 
                           B2 => n4, ZN => n11);
   U15 : INV_X1 port map( A => n11, ZN => n75);
   U16 : AOI22_X1 port map( A1 => DATA_OUT_1_port, A2 => n7, B1 => DATA_IN(1), 
                           B2 => n4, ZN => n12);
   U17 : INV_X1 port map( A => n12, ZN => n74);
   U18 : AOI22_X1 port map( A1 => DATA_OUT_2_port, A2 => n7, B1 => DATA_IN(2), 
                           B2 => n4, ZN => n13);
   U19 : INV_X1 port map( A => n13, ZN => n73);
   U20 : AOI22_X1 port map( A1 => DATA_OUT_3_port, A2 => n7, B1 => DATA_IN(3), 
                           B2 => n4, ZN => n14);
   U21 : INV_X1 port map( A => n14, ZN => n72);
   U22 : AOI22_X1 port map( A1 => DATA_OUT_4_port, A2 => n7, B1 => DATA_IN(4), 
                           B2 => n4, ZN => n15);
   U23 : INV_X1 port map( A => n15, ZN => n71);
   U24 : AOI22_X1 port map( A1 => DATA_OUT_5_port, A2 => n7, B1 => DATA_IN(5), 
                           B2 => n4, ZN => n16);
   U25 : INV_X1 port map( A => n16, ZN => n70);
   U26 : AOI22_X1 port map( A1 => DATA_OUT_6_port, A2 => n7, B1 => DATA_IN(6), 
                           B2 => n4, ZN => n17);
   U27 : INV_X1 port map( A => n17, ZN => n69);
   U28 : AOI22_X1 port map( A1 => DATA_OUT_7_port, A2 => n7, B1 => DATA_IN(7), 
                           B2 => n4, ZN => n18);
   U29 : INV_X1 port map( A => n18, ZN => n68);
   U30 : AOI22_X1 port map( A1 => DATA_OUT_8_port, A2 => n7, B1 => DATA_IN(8), 
                           B2 => n4, ZN => n19);
   U31 : INV_X1 port map( A => n19, ZN => n67);
   U32 : AOI22_X1 port map( A1 => DATA_OUT_9_port, A2 => n7, B1 => DATA_IN(9), 
                           B2 => n4, ZN => n20);
   U33 : INV_X1 port map( A => n20, ZN => n66);
   U34 : AOI22_X1 port map( A1 => DATA_OUT_10_port, A2 => n7, B1 => DATA_IN(10)
                           , B2 => n4, ZN => n21);
   U35 : INV_X1 port map( A => n21, ZN => n65);
   U36 : AOI22_X1 port map( A1 => DATA_OUT_11_port, A2 => n7, B1 => DATA_IN(11)
                           , B2 => n4, ZN => n22);
   U37 : INV_X1 port map( A => n22, ZN => n64);
   U38 : AOI22_X1 port map( A1 => DATA_OUT_12_port, A2 => n8, B1 => DATA_IN(12)
                           , B2 => n5, ZN => n23);
   U39 : INV_X1 port map( A => n23, ZN => n63);
   U40 : AOI22_X1 port map( A1 => DATA_OUT_13_port, A2 => n8, B1 => DATA_IN(13)
                           , B2 => n5, ZN => n24);
   U41 : INV_X1 port map( A => n24, ZN => n62);
   U42 : AOI22_X1 port map( A1 => DATA_OUT_14_port, A2 => n8, B1 => DATA_IN(14)
                           , B2 => n5, ZN => n25);
   U43 : INV_X1 port map( A => n25, ZN => n61);
   U44 : AOI22_X1 port map( A1 => DATA_OUT_15_port, A2 => n8, B1 => DATA_IN(15)
                           , B2 => n5, ZN => n26);
   U45 : INV_X1 port map( A => n26, ZN => n60);
   U46 : AOI22_X1 port map( A1 => DATA_OUT_16_port, A2 => n8, B1 => DATA_IN(16)
                           , B2 => n5, ZN => n27);
   U47 : INV_X1 port map( A => n27, ZN => n59);
   U48 : AOI22_X1 port map( A1 => DATA_OUT_17_port, A2 => n8, B1 => DATA_IN(17)
                           , B2 => n5, ZN => n28);
   U49 : INV_X1 port map( A => n28, ZN => n58);
   U50 : AOI22_X1 port map( A1 => DATA_OUT_18_port, A2 => n8, B1 => DATA_IN(18)
                           , B2 => n5, ZN => n29);
   U51 : INV_X1 port map( A => n29, ZN => n57);
   U52 : AOI22_X1 port map( A1 => DATA_OUT_19_port, A2 => n8, B1 => DATA_IN(19)
                           , B2 => n5, ZN => n30);
   U53 : INV_X1 port map( A => n30, ZN => n56);
   U54 : AOI22_X1 port map( A1 => DATA_OUT_20_port, A2 => n8, B1 => DATA_IN(20)
                           , B2 => n5, ZN => n31);
   U55 : INV_X1 port map( A => n31, ZN => n55);
   U56 : AOI22_X1 port map( A1 => DATA_OUT_21_port, A2 => n8, B1 => DATA_IN(21)
                           , B2 => n5, ZN => n32);
   U57 : INV_X1 port map( A => n32, ZN => n54);
   U58 : AOI22_X1 port map( A1 => DATA_OUT_22_port, A2 => n8, B1 => DATA_IN(22)
                           , B2 => n5, ZN => n33);
   U59 : INV_X1 port map( A => n33, ZN => n53);
   U60 : AOI22_X1 port map( A1 => DATA_OUT_23_port, A2 => n8, B1 => DATA_IN(23)
                           , B2 => n5, ZN => n34);
   U61 : INV_X1 port map( A => n34, ZN => n52);
   U62 : AOI22_X1 port map( A1 => DATA_OUT_24_port, A2 => n9, B1 => DATA_IN(24)
                           , B2 => n6, ZN => n35);
   U63 : INV_X1 port map( A => n35, ZN => n51);
   U64 : AOI22_X1 port map( A1 => DATA_OUT_25_port, A2 => n9, B1 => DATA_IN(25)
                           , B2 => n6, ZN => n36);
   U65 : INV_X1 port map( A => n36, ZN => n50);
   U66 : AOI22_X1 port map( A1 => DATA_OUT_26_port, A2 => n9, B1 => DATA_IN(26)
                           , B2 => n6, ZN => n37);
   U67 : INV_X1 port map( A => n37, ZN => n49);
   U68 : AOI22_X1 port map( A1 => DATA_OUT_27_port, A2 => n9, B1 => DATA_IN(27)
                           , B2 => n6, ZN => n38);
   U69 : INV_X1 port map( A => n38, ZN => n48);
   U70 : AOI22_X1 port map( A1 => DATA_OUT_28_port, A2 => n9, B1 => DATA_IN(28)
                           , B2 => n6, ZN => n39);
   U71 : INV_X1 port map( A => n39, ZN => n47);
   U72 : AOI22_X1 port map( A1 => DATA_OUT_29_port, A2 => n9, B1 => DATA_IN(29)
                           , B2 => n6, ZN => n40);
   U73 : INV_X1 port map( A => n40, ZN => n46);
   U74 : AOI22_X1 port map( A1 => DATA_OUT_30_port, A2 => n9, B1 => DATA_IN(30)
                           , B2 => n6, ZN => n41);
   U75 : INV_X1 port map( A => n41, ZN => n45);
   U76 : AOI22_X1 port map( A1 => DATA_OUT_31_port, A2 => n9, B1 => DATA_IN(31)
                           , B2 => n6, ZN => n43);
   U77 : INV_X1 port map( A => n43, ZN => n44);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_4 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_4;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, 
      n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, 
      n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, 
      n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100 : 
      std_logic;

begin
   DATA_OUT <= ( DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port );
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n44, CK => CLK, Q => 
                           DATA_OUT_31_port, QN => n_1069);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n45, CK => CLK, Q => 
                           DATA_OUT_30_port, QN => n_1070);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n46, CK => CLK, Q => 
                           DATA_OUT_29_port, QN => n_1071);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n47, CK => CLK, Q => 
                           DATA_OUT_28_port, QN => n_1072);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n48, CK => CLK, Q => 
                           DATA_OUT_27_port, QN => n_1073);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n49, CK => CLK, Q => 
                           DATA_OUT_26_port, QN => n_1074);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n50, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_1075);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n51, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n_1076);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n52, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_1077);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n53, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n_1078);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n54, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n_1079);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n55, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_1080);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n56, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_1081);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n57, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_1082);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n58, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_1083);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n59, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n_1084);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n60, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n_1085);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n61, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n_1086);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n62, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n_1087);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n63, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n_1088);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n64, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n_1089);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n65, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n_1090);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n66, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n_1091);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n67, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n_1092);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n_1093);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n_1094);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT_5_port, QN => n_1095);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_1096);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_1097);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_1098);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_1099);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_1100);
   U3 : BUF_X2 port map( A => n42, Z => n7);
   U4 : BUF_X2 port map( A => n42, Z => n8);
   U5 : BUF_X1 port map( A => n1, Z => n4);
   U6 : BUF_X1 port map( A => n1, Z => n5);
   U7 : BUF_X1 port map( A => n42, Z => n9);
   U8 : BUF_X1 port map( A => n1, Z => n6);
   U9 : AND2_X1 port map( A1 => n2, A2 => n10, ZN => n1);
   U10 : INV_X1 port map( A => n3, ZN => n2);
   U11 : INV_X1 port map( A => RST, ZN => n3);
   U12 : OR2_X1 port map( A1 => EN, A2 => n3, ZN => n10);
   U13 : INV_X1 port map( A => n10, ZN => n42);
   U14 : AOI22_X1 port map( A1 => DATA_OUT_0_port, A2 => n7, B1 => DATA_IN(0), 
                           B2 => n4, ZN => n11);
   U15 : INV_X1 port map( A => n11, ZN => n75);
   U16 : AOI22_X1 port map( A1 => DATA_OUT_1_port, A2 => n7, B1 => DATA_IN(1), 
                           B2 => n4, ZN => n12);
   U17 : INV_X1 port map( A => n12, ZN => n74);
   U18 : AOI22_X1 port map( A1 => DATA_OUT_2_port, A2 => n7, B1 => DATA_IN(2), 
                           B2 => n4, ZN => n13);
   U19 : INV_X1 port map( A => n13, ZN => n73);
   U20 : AOI22_X1 port map( A1 => DATA_OUT_3_port, A2 => n7, B1 => DATA_IN(3), 
                           B2 => n4, ZN => n14);
   U21 : INV_X1 port map( A => n14, ZN => n72);
   U22 : AOI22_X1 port map( A1 => DATA_OUT_4_port, A2 => n7, B1 => DATA_IN(4), 
                           B2 => n4, ZN => n15);
   U23 : INV_X1 port map( A => n15, ZN => n71);
   U24 : AOI22_X1 port map( A1 => DATA_OUT_5_port, A2 => n7, B1 => DATA_IN(5), 
                           B2 => n4, ZN => n16);
   U25 : INV_X1 port map( A => n16, ZN => n70);
   U26 : AOI22_X1 port map( A1 => DATA_OUT_6_port, A2 => n7, B1 => DATA_IN(6), 
                           B2 => n4, ZN => n17);
   U27 : INV_X1 port map( A => n17, ZN => n69);
   U28 : AOI22_X1 port map( A1 => DATA_OUT_7_port, A2 => n7, B1 => DATA_IN(7), 
                           B2 => n4, ZN => n18);
   U29 : INV_X1 port map( A => n18, ZN => n68);
   U30 : AOI22_X1 port map( A1 => DATA_OUT_8_port, A2 => n7, B1 => DATA_IN(8), 
                           B2 => n4, ZN => n19);
   U31 : INV_X1 port map( A => n19, ZN => n67);
   U32 : AOI22_X1 port map( A1 => DATA_OUT_9_port, A2 => n7, B1 => DATA_IN(9), 
                           B2 => n4, ZN => n20);
   U33 : INV_X1 port map( A => n20, ZN => n66);
   U34 : AOI22_X1 port map( A1 => DATA_OUT_10_port, A2 => n7, B1 => DATA_IN(10)
                           , B2 => n4, ZN => n21);
   U35 : INV_X1 port map( A => n21, ZN => n65);
   U36 : AOI22_X1 port map( A1 => DATA_OUT_11_port, A2 => n7, B1 => DATA_IN(11)
                           , B2 => n4, ZN => n22);
   U37 : INV_X1 port map( A => n22, ZN => n64);
   U38 : AOI22_X1 port map( A1 => DATA_OUT_12_port, A2 => n8, B1 => DATA_IN(12)
                           , B2 => n5, ZN => n23);
   U39 : INV_X1 port map( A => n23, ZN => n63);
   U40 : AOI22_X1 port map( A1 => DATA_OUT_13_port, A2 => n8, B1 => DATA_IN(13)
                           , B2 => n5, ZN => n24);
   U41 : INV_X1 port map( A => n24, ZN => n62);
   U42 : AOI22_X1 port map( A1 => DATA_OUT_14_port, A2 => n8, B1 => DATA_IN(14)
                           , B2 => n5, ZN => n25);
   U43 : INV_X1 port map( A => n25, ZN => n61);
   U44 : AOI22_X1 port map( A1 => DATA_OUT_15_port, A2 => n8, B1 => DATA_IN(15)
                           , B2 => n5, ZN => n26);
   U45 : INV_X1 port map( A => n26, ZN => n60);
   U46 : AOI22_X1 port map( A1 => DATA_OUT_16_port, A2 => n8, B1 => DATA_IN(16)
                           , B2 => n5, ZN => n27);
   U47 : INV_X1 port map( A => n27, ZN => n59);
   U48 : AOI22_X1 port map( A1 => DATA_OUT_17_port, A2 => n8, B1 => DATA_IN(17)
                           , B2 => n5, ZN => n28);
   U49 : INV_X1 port map( A => n28, ZN => n58);
   U50 : AOI22_X1 port map( A1 => DATA_OUT_18_port, A2 => n8, B1 => DATA_IN(18)
                           , B2 => n5, ZN => n29);
   U51 : INV_X1 port map( A => n29, ZN => n57);
   U52 : AOI22_X1 port map( A1 => DATA_OUT_19_port, A2 => n8, B1 => DATA_IN(19)
                           , B2 => n5, ZN => n30);
   U53 : INV_X1 port map( A => n30, ZN => n56);
   U54 : AOI22_X1 port map( A1 => DATA_OUT_20_port, A2 => n8, B1 => DATA_IN(20)
                           , B2 => n5, ZN => n31);
   U55 : INV_X1 port map( A => n31, ZN => n55);
   U56 : AOI22_X1 port map( A1 => DATA_OUT_21_port, A2 => n8, B1 => DATA_IN(21)
                           , B2 => n5, ZN => n32);
   U57 : INV_X1 port map( A => n32, ZN => n54);
   U58 : AOI22_X1 port map( A1 => DATA_OUT_22_port, A2 => n8, B1 => DATA_IN(22)
                           , B2 => n5, ZN => n33);
   U59 : INV_X1 port map( A => n33, ZN => n53);
   U60 : AOI22_X1 port map( A1 => DATA_OUT_23_port, A2 => n8, B1 => DATA_IN(23)
                           , B2 => n5, ZN => n34);
   U61 : INV_X1 port map( A => n34, ZN => n52);
   U62 : AOI22_X1 port map( A1 => DATA_OUT_24_port, A2 => n9, B1 => DATA_IN(24)
                           , B2 => n6, ZN => n35);
   U63 : INV_X1 port map( A => n35, ZN => n51);
   U64 : AOI22_X1 port map( A1 => DATA_OUT_25_port, A2 => n9, B1 => DATA_IN(25)
                           , B2 => n6, ZN => n36);
   U65 : INV_X1 port map( A => n36, ZN => n50);
   U66 : AOI22_X1 port map( A1 => DATA_OUT_26_port, A2 => n9, B1 => DATA_IN(26)
                           , B2 => n6, ZN => n37);
   U67 : INV_X1 port map( A => n37, ZN => n49);
   U68 : AOI22_X1 port map( A1 => DATA_OUT_27_port, A2 => n9, B1 => DATA_IN(27)
                           , B2 => n6, ZN => n38);
   U69 : INV_X1 port map( A => n38, ZN => n48);
   U70 : AOI22_X1 port map( A1 => DATA_OUT_28_port, A2 => n9, B1 => DATA_IN(28)
                           , B2 => n6, ZN => n39);
   U71 : INV_X1 port map( A => n39, ZN => n47);
   U72 : AOI22_X1 port map( A1 => DATA_OUT_29_port, A2 => n9, B1 => DATA_IN(29)
                           , B2 => n6, ZN => n40);
   U73 : INV_X1 port map( A => n40, ZN => n46);
   U74 : AOI22_X1 port map( A1 => DATA_OUT_30_port, A2 => n9, B1 => DATA_IN(30)
                           , B2 => n6, ZN => n41);
   U75 : INV_X1 port map( A => n41, ZN => n45);
   U76 : AOI22_X1 port map( A1 => DATA_OUT_31_port, A2 => n9, B1 => DATA_IN(31)
                           , B2 => n6, ZN => n43);
   U77 : INV_X1 port map( A => n43, ZN => n44);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_cmp6_3 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end ALU_N32_DW01_cmp6_3;

architecture SYN_rpl of ALU_N32_DW01_cmp6_3 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44 : 
      std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B(24), B => A(24), ZN => n27);
   U2 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n37);
   U3 : XNOR2_X1 port map( A => B(23), B => A(23), ZN => n28);
   U4 : XNOR2_X1 port map( A => B(21), B => A(21), ZN => n30);
   U5 : XNOR2_X1 port map( A => B(20), B => A(20), ZN => n31);
   U6 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n10);
   U7 : XNOR2_X1 port map( A => B(28), B => A(28), ZN => n41);
   U8 : XNOR2_X1 port map( A => B(29), B => A(29), ZN => n40);
   U9 : XNOR2_X1 port map( A => B(17), B => A(17), ZN => n34);
   U10 : XNOR2_X1 port map( A => B(16), B => A(16), ZN => n17);
   U11 : XNOR2_X1 port map( A => B(30), B => A(30), ZN => n38);
   U12 : XNOR2_X1 port map( A => B(27), B => A(27), ZN => n42);
   U13 : XNOR2_X1 port map( A => B(26), B => A(26), ZN => n43);
   U14 : XNOR2_X1 port map( A => B(9), B => A(9), ZN => n23);
   U15 : XNOR2_X1 port map( A => B(11), B => A(11), ZN => n22);
   U16 : XNOR2_X1 port map( A => B(19), B => A(19), ZN => n32);
   U17 : XNOR2_X1 port map( A => B(25), B => A(25), ZN => n44);
   U18 : XNOR2_X1 port map( A => B(10), B => A(10), ZN => n39);
   U19 : XNOR2_X1 port map( A => B(18), B => A(18), ZN => n33);
   U20 : XNOR2_X1 port map( A => B(13), B => A(13), ZN => n20);
   U21 : XNOR2_X1 port map( A => B(15), B => A(15), ZN => n18);
   U22 : XNOR2_X1 port map( A => B(22), B => A(22), ZN => n29);
   U23 : XNOR2_X1 port map( A => B(7), B => A(7), ZN => n7);
   U24 : XNOR2_X1 port map( A => B(12), B => A(12), ZN => n21);
   U25 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n9);
   U26 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n11);
   U27 : XNOR2_X1 port map( A => B(14), B => A(14), ZN => n19);
   U28 : XNOR2_X1 port map( A => B(0), B => A(0), ZN => n14);
   U29 : XNOR2_X1 port map( A => B(8), B => A(8), ZN => n24);
   U30 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n13);
   U31 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n8);
   U32 : XNOR2_X1 port map( A => B(1), B => A(1), ZN => n12);
   U33 : NAND4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => NE);
   U34 : NOR2_X1 port map( A1 => n5, A2 => n6, ZN => n4);
   U35 : NAND4_X1 port map( A1 => n7, A2 => n8, A3 => n9, A4 => n10, ZN => n6);
   U36 : NAND4_X1 port map( A1 => n11, A2 => n12, A3 => n13, A4 => n14, ZN => 
                           n5);
   U37 : NOR2_X1 port map( A1 => n15, A2 => n16, ZN => n3);
   U38 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           n16);
   U39 : NAND4_X1 port map( A1 => n21, A2 => n22, A3 => n23, A4 => n24, ZN => 
                           n15);
   U40 : NOR2_X1 port map( A1 => n25, A2 => n26, ZN => n2);
   U41 : NAND4_X1 port map( A1 => n27, A2 => n28, A3 => n29, A4 => n30, ZN => 
                           n26);
   U42 : NAND4_X1 port map( A1 => n31, A2 => n32, A3 => n33, A4 => n34, ZN => 
                           n25);
   U43 : NOR2_X1 port map( A1 => n35, A2 => n36, ZN => n1);
   U44 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           n36);
   U45 : NAND4_X1 port map( A1 => n41, A2 => n42, A3 => n43, A4 => n44, ZN => 
                           n35);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_cmp6_2 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end ALU_N32_DW01_cmp6_2;

architecture SYN_rpl of ALU_N32_DW01_cmp6_2 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437 : 
      std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => n158);
   U2 : NAND2_X1 port map( A1 => n420, A2 => n182, ZN => n415);
   U3 : INV_X1 port map( A => n11, ZN => n42);
   U4 : AND2_X1 port map( A1 => n121, A2 => n122, ZN => n1);
   U5 : XOR2_X1 port map( A => B(31), B => A(31), Z => n2);
   U6 : AND2_X1 port map( A1 => A(17), A2 => n355, ZN => n3);
   U7 : NAND2_X1 port map( A1 => n98, A2 => n286, ZN => n33);
   U8 : OR2_X1 port map( A1 => n298, A2 => n222, ZN => n4);
   U9 : OR2_X1 port map( A1 => n229, A2 => n33, ZN => n5);
   U10 : AND2_X1 port map( A1 => B(9), A2 => n434, ZN => n6);
   U11 : NAND2_X1 port map( A1 => n121, A2 => n122, ZN => n7);
   U12 : AND3_X1 port map( A1 => n417, A2 => n181, A3 => n213, ZN => n8);
   U13 : INV_X1 port map( A => n36, ZN => n9);
   U14 : INV_X2 port map( A => n9, ZN => n10);
   U15 : NAND2_X1 port map( A1 => B(25), A2 => n427, ZN => n36);
   U16 : AND4_X2 port map( A1 => n132, A2 => n133, A3 => n134, A4 => n135, ZN 
                           => n11);
   U17 : INV_X1 port map( A => n55, ZN => n12);
   U18 : INV_X1 port map( A => n55, ZN => n13);
   U19 : NAND2_X2 port map( A1 => n128, A2 => n307, ZN => n55);
   U20 : AND2_X2 port map( A1 => n98, A2 => n286, ZN => n14);
   U21 : OAI211_X1 port map( C1 => n361, C2 => n362, A => n245, B => n66, ZN =>
                           n222);
   U22 : NOR2_X1 port map( A1 => n297, A2 => n4, ZN => n296);
   U23 : INV_X2 port map( A => n228, ZN => n121);
   U24 : NAND2_X2 port map( A1 => n60, A2 => n253, ZN => n67);
   U25 : NAND2_X2 port map( A1 => n424, A2 => n178, ZN => n226);
   U26 : AND2_X1 port map( A1 => n188, A2 => n15, ZN => n184);
   U27 : AND2_X1 port map( A1 => n146, A2 => n152, ZN => n15);
   U28 : AND2_X1 port map( A1 => n16, A2 => n151, ZN => n189);
   U29 : OR2_X1 port map( A1 => n211, A2 => n212, ZN => n16);
   U30 : OR2_X1 port map( A1 => B(31), A2 => n131, ZN => n35);
   U31 : NAND2_X1 port map( A1 => n121, A2 => n122, ZN => n32);
   U32 : NOR2_X1 port map( A1 => n222, A2 => n287, ZN => n281);
   U33 : AOI21_X1 port map( B1 => n280, B2 => n281, A => n282, ZN => n279);
   U34 : AOI21_X1 port map( B1 => n108, B2 => n11, A => n109, ZN => n90);
   U35 : NOR3_X1 port map( A1 => n115, A2 => n116, A3 => n117, ZN => n108);
   U36 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => n109);
   U37 : AOI21_X1 port map( B1 => n92, B2 => n93, A => n94, ZN => n91);
   U38 : NAND2_X1 port map( A1 => n95, A2 => n96, ZN => n94);
   U39 : NOR2_X1 port map( A1 => n101, A2 => n42, ZN => n92);
   U40 : AND4_X1 port map( A1 => n99, A2 => n83, A3 => n12, A4 => n41, ZN => 
                           n93);
   U41 : AOI22_X1 port map( A1 => n76, A2 => n77, B1 => n78, B2 => n79, ZN => 
                           n23);
   U42 : NOR2_X1 port map( A1 => n84, A2 => n85, ZN => n77);
   U43 : NOR2_X1 port map( A1 => n80, A2 => n81, ZN => n79);
   U44 : NOR2_X1 port map( A1 => n86, A2 => n42, ZN => n76);
   U45 : NOR2_X1 port map( A1 => n170, A2 => n149, ZN => n192);
   U46 : NOR2_X1 port map( A1 => n263, A2 => n224, ZN => n262);
   U47 : NOR2_X1 port map( A1 => n222, A2 => n271, ZN => n270);
   U48 : NOR2_X1 port map( A1 => n222, A2 => n224, ZN => n315);
   U49 : NOR2_X1 port map( A1 => n67, A2 => n229, ZN => n293);
   U50 : AOI21_X1 port map( B1 => n141, B2 => n142, A => n143, ZN => n125);
   U51 : NOR2_X1 port map( A1 => n153, A2 => n154, ZN => n124);
   U52 : NOR2_X1 port map( A1 => n42, A2 => n127, ZN => n126);
   U53 : AOI21_X1 port map( B1 => n398, B2 => n399, A => n400, ZN => n367);
   U54 : NOR2_X1 port map( A1 => n326, A2 => n412, ZN => n398);
   U55 : NOR2_X1 port map( A1 => n407, A2 => n408, ZN => n399);
   U56 : NOR2_X1 port map( A1 => n326, A2 => n401, ZN => n400);
   U57 : NOR2_X1 port map( A1 => n267, A2 => n106, ZN => n294);
   U58 : NOR2_X1 port map( A1 => n55, A2 => n222, ZN => n221);
   U59 : OAI211_X1 port map( C1 => n88, C2 => n89, A => n90, B => n91, ZN => 
                           n21);
   U60 : NAND4_X1 port map( A1 => n50, A2 => n51, A3 => n52, A4 => n53, ZN => 
                           n24);
   U61 : NOR2_X1 port map( A1 => n364, A2 => n59, ZN => n58);
   U62 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => n56);
   U63 : AOI21_X1 port map( B1 => n63, B2 => n64, A => n65, ZN => n57);
   U64 : NAND2_X1 port map( A1 => n248, A2 => n226, ZN => n247);
   U65 : NAND2_X1 port map( A1 => n304, A2 => n226, ZN => n302);
   U66 : NOR2_X1 port map( A1 => n267, A2 => n106, ZN => n304);
   U67 : NOR2_X1 port map( A1 => n295, A2 => n296, ZN => n278);
   U68 : NOR3_X1 port map( A1 => n305, A2 => n222, A3 => n306, ZN => n295);
   U69 : NOR2_X1 port map( A1 => n318, A2 => n319, ZN => n317);
   U70 : OAI21_X1 port map( B1 => n326, B2 => n329, A => n330, ZN => n318);
   U71 : NAND2_X1 port map( A1 => n320, A2 => n321, ZN => n319);
   U72 : NOR2_X1 port map( A1 => n331, A2 => n67, ZN => n330);
   U73 : INV_X1 port map( A => n67, ZN => n64);
   U74 : INV_X1 port map( A => n67, ZN => n72);
   U75 : NOR2_X1 port map( A1 => n130, A2 => n5, ZN => n316);
   U76 : INV_X1 port map( A => n170, ZN => n185);
   U77 : INV_X1 port map( A => n122, ZN => n143);
   U78 : INV_X1 port map( A => n149, ZN => n159);
   U79 : AND2_X1 port map( A1 => n37, A2 => n44, ZN => n176);
   U80 : NOR2_X1 port map( A1 => n138, A2 => n139, ZN => n132);
   U81 : NAND2_X1 port map( A1 => n180, A2 => n193, ZN => n149);
   U82 : NAND2_X1 port map( A1 => n353, A2 => n354, ZN => n224);
   U83 : NOR2_X1 port map( A1 => n249, A2 => n357, ZN => n353);
   U84 : AND2_X1 port map( A1 => n61, A2 => n66, ZN => n177);
   U85 : NAND2_X1 port map( A1 => n273, A2 => n34, ZN => n106);
   U86 : NAND2_X1 port map( A1 => n259, A2 => n69, ZN => n229);
   U87 : NOR3_X1 port map( A1 => n250, A2 => n251, A3 => n252, ZN => n246);
   U88 : OAI21_X1 port map( B1 => n67, B2 => n257, A => n10, ZN => n250);
   U89 : NOR2_X1 port map( A1 => n67, A2 => n70, ZN => n251);
   U90 : NOR3_X1 port map( A1 => n223, A2 => n224, A3 => n140, ZN => n220);
   U91 : NOR2_X1 port map( A1 => n229, A2 => n67, ZN => n225);
   U92 : NOR2_X1 port map( A1 => n33, A2 => n228, ZN => n227);
   U93 : NOR3_X1 port map( A1 => n272, A2 => n224, A3 => n273, ZN => n269);
   U94 : NOR2_X1 port map( A1 => n267, A2 => n67, ZN => n274);
   U95 : NOR2_X1 port map( A1 => n229, A2 => n33, ZN => n275);
   U96 : NOR2_X1 port map( A1 => n375, A2 => n326, ZN => n370);
   U97 : NOR3_X1 port map( A1 => n26, A2 => n27, A3 => n28, ZN => n25);
   U98 : OAI21_X1 port map( B1 => n45, B2 => n46, A => n47, ZN => n26);
   U99 : NOR2_X1 port map( A1 => n38, A2 => n39, ZN => n27);
   U100 : NOR2_X1 port map( A1 => n29, A2 => n30, ZN => n28);
   U101 : NAND4_X1 port map( A1 => n31, A2 => n119, A3 => n41, A4 => n11, ZN =>
                           n30);
   U102 : NOR2_X1 port map( A1 => n33, A2 => n34, ZN => n31);
   U103 : NAND4_X1 port map( A1 => n40, A2 => n13, A3 => n41, A4 => n11, ZN => 
                           n39);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n43, ZN => n40);
   U105 : INV_X1 port map( A => n7, ZN => n41);
   U106 : INV_X1 port map( A => n181, ZN => n179);
   U107 : OAI21_X1 port map( B1 => n155, B2 => n156, A => n157, ZN => n154);
   U108 : NAND4_X1 port map( A1 => n147, A2 => n146, A3 => n159, A4 => n6, ZN 
                           => n157);
   U109 : NAND4_X1 port map( A1 => n44, A2 => n10, A3 => n35, A4 => n37, ZN => 
                           n38);
   U110 : NAND4_X1 port map( A1 => n128, A2 => n14, A3 => n35, A4 => n129, ZN 
                           => n127);
   U111 : INV_X1 port map( A => n130, ZN => n129);
   U112 : NAND2_X1 port map( A1 => n417, A2 => n147, ZN => n182);
   U113 : NOR2_X1 port map( A1 => n82, A2 => n42, ZN => n78);
   U114 : NAND4_X1 port map( A1 => n3, A2 => n83, A3 => n119, A4 => n1, ZN => 
                           n82);
   U115 : INV_X1 port map( A => n33, ZN => n83);
   U116 : NAND4_X1 port map( A1 => n74, A2 => n349, A3 => n119, A4 => n113, ZN 
                           => n110);
   U117 : INV_X1 port map( A => n45, ZN => n113);
   U118 : NOR2_X1 port map( A1 => n222, A2 => n264, ZN => n261);
   U119 : NAND4_X1 port map( A1 => n265, A2 => n134, A3 => n266, A4 => n226, ZN
                           => n264);
   U120 : NOR2_X1 port map( A1 => n137, A2 => n229, ZN => n265);
   U121 : NOR2_X1 port map( A1 => n267, A2 => n106, ZN => n266);
   U122 : NAND2_X1 port map( A1 => n292, A2 => n43, ZN => n105);
   U123 : OAI211_X1 port map( C1 => n202, C2 => n393, A => n158, B => n394, ZN 
                           => n381);
   U124 : NAND2_X1 port map( A1 => n199, A2 => n200, ZN => n393);
   U125 : NAND4_X1 port map( A1 => n102, A2 => n44, A3 => n37, A4 => n103, ZN 
                           => n101);
   U126 : AND2_X1 port map( A1 => n10, A2 => n107, ZN => n102);
   U127 : NOR2_X1 port map( A1 => n104, A2 => n105, ZN => n103);
   U128 : NOR2_X1 port map( A1 => n149, A2 => n150, ZN => n141);
   U129 : NAND2_X1 port map( A1 => n151, A2 => n152, ZN => n150);
   U130 : AOI21_X1 port map( B1 => n230, B2 => n231, A => n232, ZN => n218);
   U131 : NOR2_X1 port map( A1 => n222, A2 => n260, ZN => n230);
   U132 : NOR2_X1 port map( A1 => n246, A2 => n247, ZN => n231);
   U133 : NOR2_X1 port map( A1 => n233, A2 => n234, ZN => n232);
   U134 : NOR2_X1 port map( A1 => n54, A2 => n55, ZN => n53);
   U135 : NAND2_X1 port map( A1 => n35, A2 => n14, ZN => n54);
   U136 : NAND2_X1 port map( A1 => n394, A2 => n152, ZN => n148);
   U137 : NAND2_X1 port map( A1 => n61, A2 => n254, ZN => n178);
   U138 : NAND4_X1 port map( A1 => n83, A2 => n12, A3 => n120, A4 => n52, ZN =>
                           n115);
   U139 : INV_X1 port map( A => n123, ZN => n120);
   U140 : INV_X1 port map( A => n55, ZN => n119);
   U141 : NOR2_X1 port map( A1 => n171, A2 => n149, ZN => n168);
   U142 : NOR2_X1 port map( A1 => n196, A2 => n197, ZN => n191);
   U143 : OAI21_X1 port map( B1 => n198, B2 => n199, A => n152, ZN => n197);
   U144 : NOR2_X1 port map( A1 => n172, A2 => n173, ZN => n166);
   U145 : NAND2_X1 port map( A1 => n183, A2 => n10, ZN => n172);
   U146 : NAND2_X1 port map( A1 => n244, A2 => n114, ZN => n228);
   U147 : AND2_X1 port map( A1 => n148, A2 => n17, ZN => n142);
   U148 : AND2_X1 port map( A1 => n146, A2 => n147, ZN => n17);
   U149 : NAND4_X1 port map( A1 => n164, A2 => n165, A3 => n166, A4 => n167, ZN
                           => n88);
   U150 : AND2_X1 port map( A1 => n107, A2 => n213, ZN => n164);
   U151 : NAND4_X1 port map( A1 => n168, A2 => n185, A3 => n169, A4 => n146, ZN
                           => n167);
   U152 : NAND4_X1 port map( A1 => n189, A2 => n190, A3 => n191, A4 => n192, ZN
                           => n165);
   U153 : NOR2_X1 port map( A1 => n6, A2 => n201, ZN => n402);
   U154 : NOR2_X1 port map( A1 => n161, A2 => n162, ZN => n153);
   U155 : NAND2_X1 port map( A1 => n163, A2 => n146, ZN => n161);
   U156 : NAND2_X1 port map( A1 => n147, A2 => n159, ZN => n162);
   U157 : NOR2_X1 port map( A1 => n68, A2 => n69, ZN => n63);
   U158 : INV_X1 port map( A => n70, ZN => n68);
   U159 : NOR2_X1 port map( A1 => n288, A2 => n289, ZN => n280);
   U160 : NAND4_X1 port map( A1 => n293, A2 => n14, A3 => n294, A4 => n226, ZN 
                           => n288);
   U161 : NAND2_X1 port map( A1 => n44, A2 => n10, ZN => n81);
   U162 : NAND2_X1 port map( A1 => n35, A2 => n10, ZN => n84);
   U163 : NAND2_X1 port map( A1 => n323, A2 => n146, ZN => n163);
   U164 : NAND2_X1 port map( A1 => n206, A2 => n207, ZN => n212);
   U165 : NAND2_X1 port map( A1 => n35, A2 => n2, ZN => n96);
   U166 : NAND2_X1 port map( A1 => n35, A2 => n118, ZN => n117);
   U167 : NAND2_X1 port map( A1 => n97, A2 => n35, ZN => n95);
   U168 : INV_X1 port map( A => n98, ZN => n97);
   U169 : NAND2_X1 port map( A1 => n35, A2 => n37, ZN => n80);
   U170 : NAND2_X1 port map( A1 => n158, A2 => n394, ZN => n412);
   U171 : NAND2_X1 port map( A1 => n386, A2 => n195, ZN => n188);
   U172 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => n59);
   U173 : NAND2_X1 port map( A1 => n112, A2 => n73, ZN => n357);
   U174 : NOR2_X1 port map( A1 => n187, A2 => n149, ZN => n186);
   U175 : NOR2_X1 port map( A1 => n107, A2 => n224, ZN => n300);
   U176 : NOR2_X1 port map( A1 => n302, A2 => n303, ZN => n299);
   U177 : NOR2_X1 port map( A1 => n310, A2 => n224, ZN => n309);
   U178 : NOR2_X1 port map( A1 => n311, A2 => n312, ZN => n308);
   U179 : NAND2_X1 port map( A1 => n342, A2 => n343, ZN => n130);
   U180 : NOR2_X1 port map( A1 => n344, A2 => n345, ZN => n343);
   U181 : NOR2_X1 port map( A1 => n349, A2 => n105, ZN => n342);
   U182 : NAND2_X1 port map( A1 => n100, A2 => n310, ZN => n345);
   U183 : NOR2_X1 port map( A1 => n327, A2 => n151, ZN => n325);
   U184 : NAND2_X1 port map( A1 => n313, A2 => n226, ZN => n311);
   U185 : NOR2_X1 port map( A1 => n106, A2 => n314, ZN => n313);
   U186 : NAND2_X1 port map( A1 => n87, A2 => n123, ZN => n314);
   U187 : NAND2_X1 port map( A1 => n323, A2 => n160, ZN => n408);
   U188 : NAND2_X1 port map( A1 => n75, A2 => n74, ZN => n139);
   U189 : INV_X1 port map( A => n35, ZN => n104);
   U190 : NOR2_X1 port map( A1 => n413, A2 => n414, ZN => n366);
   U191 : NOR2_X1 port map( A1 => n326, A2 => n429, ZN => n413);
   U192 : NAND4_X1 port map( A1 => n226, A2 => n44, A3 => n415, A4 => n416, ZN 
                           => n414);
   U193 : NOR2_X1 port map( A1 => n243, A2 => n244, ZN => n242);
   U194 : OR3_X1 port map( A1 => n112, A2 => n55, A3 => n45, ZN => n111);
   U195 : NAND2_X1 port map( A1 => n70, A2 => n140, ZN => n138);
   U196 : NAND4_X1 port map( A1 => n267, A2 => n83, A3 => n13, A4 => n1, ZN => 
                           n86);
   U197 : INV_X1 port map( A => n66, ZN => n65);
   U198 : NAND2_X1 port map( A1 => n322, A2 => n8, ZN => n321);
   U199 : AND2_X1 port map( A1 => n163, A2 => n323, ZN => n322);
   U200 : NAND2_X1 port map( A1 => n188, A2 => n386, ZN => n407);
   U201 : AND2_X1 port map( A1 => n417, A2 => n213, ZN => n420);
   U202 : INV_X1 port map( A => n73, ZN => n71);
   U203 : NAND2_X1 port map( A1 => n334, A2 => n335, ZN => n329);
   U204 : NOR2_X1 port map( A1 => n327, A2 => n194, ZN => n335);
   U205 : OR2_X1 port map( A1 => n48, A2 => n45, ZN => n47);
   U206 : AND2_X1 port map( A1 => n151, A2 => n152, ZN => n169);
   U207 : NAND2_X1 port map( A1 => n283, A2 => n284, ZN => n282);
   U208 : NAND2_X1 port map( A1 => n285, A2 => n245, ZN => n283);
   U209 : NAND2_X1 port map( A1 => n245, A2 => n2, ZN => n284);
   U210 : AND4_X1 port map( A1 => n74, A2 => n75, A3 => n10, A4 => n37, ZN => 
                           n50);
   U211 : INV_X1 port map( A => n100, ZN => n99);
   U212 : INV_X1 port map( A => B(12), ZN => n421);
   U213 : INV_X1 port map( A => B(9), ZN => n328);
   U214 : NAND2_X1 port map( A1 => A(10), A2 => n324, ZN => n146);
   U215 : INV_X1 port map( A => B(19), ZN => n372);
   U216 : INV_X1 port map( A => B(26), ZN => n352);
   U217 : INV_X1 port map( A => B(27), ZN => n359);
   U218 : NAND2_X1 port map( A1 => A(24), A2 => n425, ZN => n61);
   U219 : INV_X1 port map( A => B(24), ZN => n425);
   U220 : INV_X1 port map( A => B(25), ZN => n363);
   U221 : INV_X1 port map( A => A(10), ZN => n431);
   U222 : NAND2_X1 port map( A1 => B(31), A2 => n131, ZN => n245);
   U223 : INV_X1 port map( A => A(31), ZN => n131);
   U224 : NAND2_X1 port map( A1 => B(27), A2 => n239, ZN => n74);
   U225 : INV_X1 port map( A => B(21), ZN => n358);
   U226 : INV_X1 port map( A => B(15), ZN => n374);
   U227 : NAND2_X1 port map( A1 => A(16), A2 => n350, ZN => n43);
   U228 : NAND2_X1 port map( A1 => B(24), A2 => n428, ZN => n254);
   U229 : INV_X1 port map( A => A(24), ZN => n428);
   U230 : INV_X1 port map( A => A(30), ZN => n338);
   U231 : NAND2_X1 port map( A1 => B(21), A2 => n256, ZN => n70);
   U232 : NAND2_X1 port map( A1 => A(23), A2 => n365, ZN => n62);
   U233 : INV_X1 port map( A => B(23), ZN => n365);
   U234 : NAND2_X1 port map( A1 => B(19), A2 => n356, ZN => n140);
   U235 : NAND2_X1 port map( A1 => B(26), A2 => n348, ZN => n244);
   U236 : INV_X1 port map( A => A(3), ZN => n391);
   U237 : INV_X1 port map( A => A(4), ZN => n389);
   U238 : NAND2_X1 port map( A1 => B(28), A2 => n238, ZN => n128);
   U239 : INV_X1 port map( A => A(17), ZN => n268);
   U240 : NAND2_X1 port map( A1 => B(14), A2 => n346, ZN => n310);
   U241 : INV_X1 port map( A => A(11), ZN => n436);
   U242 : INV_X1 port map( A => A(16), ZN => n351);
   U243 : INV_X1 port map( A => B(14), ZN => n347);
   U244 : NAND2_X1 port map( A1 => B(23), A2 => n255, ZN => n145);
   U245 : INV_X1 port map( A => A(23), ZN => n255);
   U246 : NAND2_X1 port map( A1 => A(4), A2 => n395, ZN => n200);
   U247 : NAND2_X1 port map( A1 => B(29), A2 => n241, ZN => n75);
   U248 : NAND2_X1 port map( A1 => A(3), A2 => n396, ZN => n199);
   U249 : NAND2_X1 port map( A1 => B(12), A2 => n437, ZN => n417);
   U250 : NAND4_X1 port map( A1 => n202, A2 => n203, A3 => n204, A4 => n205, ZN
                           => n190);
   U251 : AND2_X1 port map( A1 => n206, A2 => n207, ZN => n205);
   U252 : NAND2_X1 port map( A1 => n209, A2 => n210, ZN => n203);
   U253 : INV_X1 port map( A => B(28), ZN => n49);
   U254 : NOR2_X1 port map( A1 => n235, A2 => n236, ZN => n234);
   U255 : OAI21_X1 port map( B1 => n55, B2 => n74, A => n237, ZN => n236);
   U256 : NAND2_X1 port map( A1 => B(28), A2 => n238, ZN => n237);
   U257 : NOR2_X1 port map( A1 => n376, A2 => n377, ZN => n375);
   U258 : OAI21_X1 port map( B1 => n378, B2 => n379, A => n380, ZN => n377);
   U259 : NAND2_X1 port map( A1 => A(30), A2 => n339, ZN => n98);
   U260 : NAND2_X1 port map( A1 => A(11), A2 => n419, ZN => n193);
   U261 : NAND2_X1 port map( A1 => B(6), A2 => n411, ZN => n386);
   U262 : NAND2_X1 port map( A1 => B(15), A2 => n301, ZN => n107);
   U263 : INV_X1 port map( A => B(29), ZN => n360);
   U264 : NAND2_X1 port map( A1 => B(20), A2 => n341, ZN => n259);
   U265 : INV_X1 port map( A => B(20), ZN => n340);
   U266 : INV_X1 port map( A => B(18), ZN => n422);
   U267 : NAND2_X1 port map( A1 => B(18), A2 => n423, ZN => n273);
   U268 : NAND2_X1 port map( A1 => B(4), A2 => n389, ZN => n206);
   U269 : INV_X1 port map( A => B(4), ZN => n395);
   U270 : NAND2_X1 port map( A1 => A(28), A2 => n49, ZN => n46);
   U271 : NAND2_X1 port map( A1 => A(28), A2 => n49, ZN => n307);
   U272 : INV_X1 port map( A => A(28), ZN => n238);
   U273 : NAND2_X1 port map( A1 => A(29), A2 => n360, ZN => n48);
   U274 : INV_X1 port map( A => A(29), ZN => n241);
   U275 : INV_X1 port map( A => B(17), ZN => n355);
   U276 : NAND2_X1 port map( A1 => B(17), A2 => n268, ZN => n137);
   U277 : NAND2_X1 port map( A1 => B(16), A2 => n351, ZN => n292);
   U278 : INV_X1 port map( A => B(16), ZN => n350);
   U279 : INV_X1 port map( A => B(13), ZN => n373);
   U280 : NAND2_X1 port map( A1 => B(13), A2 => n435, ZN => n213);
   U281 : INV_X1 port map( A => A(21), ZN => n256);
   U282 : NAND2_X1 port map( A1 => A(21), A2 => n358, ZN => n73);
   U283 : NAND2_X1 port map( A1 => B(30), A2 => n338, ZN => n286);
   U284 : INV_X1 port map( A => B(30), ZN => n339);
   U285 : INV_X1 port map( A => A(20), ZN => n341);
   U286 : NAND2_X1 port map( A1 => A(20), A2 => n340, ZN => n69);
   U287 : NAND2_X1 port map( A1 => B(22), A2 => n332, ZN => n253);
   U288 : INV_X1 port map( A => B(22), ZN => n333);
   U289 : NAND2_X1 port map( A1 => A(27), A2 => n359, ZN => n112);
   U290 : INV_X1 port map( A => A(27), ZN => n239);
   U291 : NAND2_X1 port map( A1 => A(26), A2 => n352, ZN => n114);
   U292 : INV_X1 port map( A => A(26), ZN => n348);
   U293 : NAND2_X1 port map( A1 => B(5), A2 => n388, ZN => n171);
   U294 : INV_X1 port map( A => B(5), ZN => n406);
   U295 : NAND2_X1 port map( A1 => A(9), A2 => n328, ZN => n151);
   U296 : INV_X1 port map( A => A(9), ZN => n434);
   U297 : INV_X1 port map( A => B(7), ZN => n336);
   U298 : NAND2_X1 port map( A1 => B(7), A2 => n409, ZN => n160);
   U299 : INV_X1 port map( A => A(2), ZN => n397);
   U300 : NAND2_X1 port map( A1 => A(2), A2 => n20, ZN => n211);
   U301 : NAND2_X1 port map( A1 => B(11), A2 => n436, ZN => n181);
   U302 : INV_X1 port map( A => B(11), ZN => n419);
   U303 : NAND2_X1 port map( A1 => A(19), A2 => n372, ZN => n87);
   U304 : INV_X1 port map( A => A(19), ZN => n356);
   U305 : NAND2_X1 port map( A1 => A(8), A2 => n432, ZN => n152);
   U306 : INV_X1 port map( A => A(8), ZN => n433);
   U307 : NAND2_X1 port map( A1 => A(25), A2 => n363, ZN => n66);
   U308 : INV_X1 port map( A => A(25), ZN => n427);
   U309 : NAND2_X1 port map( A1 => B(10), A2 => n431, ZN => n323);
   U310 : INV_X1 port map( A => B(10), ZN => n324);
   U311 : NAND2_X1 port map( A1 => A(18), A2 => n422, ZN => n34);
   U312 : INV_X1 port map( A => A(18), ZN => n423);
   U313 : NAND2_X1 port map( A1 => A(13), A2 => n373, ZN => n180);
   U314 : INV_X1 port map( A => A(13), ZN => n435);
   U315 : INV_X1 port map( A => A(15), ZN => n301);
   U316 : NAND2_X1 port map( A1 => A(15), A2 => n374, ZN => n123);
   U317 : INV_X1 port map( A => B(6), ZN => n410);
   U318 : NAND2_X1 port map( A1 => A(22), A2 => n333, ZN => n60);
   U319 : INV_X1 port map( A => A(22), ZN => n332);
   U320 : INV_X1 port map( A => A(7), ZN => n409);
   U321 : NAND2_X1 port map( A1 => A(7), A2 => n336, ZN => n194);
   U322 : NAND2_X1 port map( A1 => A(12), A2 => n421, ZN => n147);
   U323 : INV_X1 port map( A => A(12), ZN => n437);
   U324 : NOR2_X1 port map( A1 => n21, A2 => n22, ZN => LE);
   U325 : NAND2_X1 port map( A1 => A(5), A2 => n406, ZN => n201);
   U326 : INV_X1 port map( A => A(5), ZN => n388);
   U327 : NAND2_X1 port map( A1 => B(3), A2 => n391, ZN => n207);
   U328 : INV_X1 port map( A => B(3), ZN => n396);
   U329 : NAND2_X1 port map( A1 => A(14), A2 => n347, ZN => n100);
   U330 : INV_X1 port map( A => A(14), ZN => n346);
   U331 : NAND2_X1 port map( A1 => A(0), A2 => n18, ZN => n210);
   U332 : NOR2_X1 port map( A1 => A(0), A2 => n18, ZN => n378);
   U333 : NAND2_X1 port map( A1 => B(8), A2 => n433, ZN => n394);
   U334 : INV_X1 port map( A => B(8), ZN => n432);
   U335 : NAND2_X1 port map( A1 => B(2), A2 => n397, ZN => n202);
   U336 : NAND2_X1 port map( A1 => A(6), A2 => n410, ZN => n195);
   U337 : INV_X1 port map( A => A(6), ZN => n411);
   U338 : NAND2_X1 port map( A1 => B(1), A2 => n208, ZN => n204);
   U339 : INV_X1 port map( A => A(1), ZN => n208);
   U340 : NAND2_X1 port map( A1 => A(1), A2 => n19, ZN => n209);
   U341 : NAND2_X1 port map( A1 => A(1), A2 => n19, ZN => n380);
   U342 : NOR2_X1 port map( A1 => A(1), A2 => n19, ZN => n379);
   U343 : INV_X1 port map( A => B(0), ZN => n18);
   U344 : INV_X1 port map( A => B(1), ZN => n19);
   U345 : INV_X1 port map( A => B(2), ZN => n20);
   U346 : NAND3_X1 port map( A1 => n23, A2 => n24, A3 => n25, ZN => n22);
   U347 : NAND3_X1 port map( A1 => n35, A2 => n10, A3 => n37, ZN => n29);
   U348 : NAND3_X1 port map( A1 => n56, A2 => n57, A3 => n58, ZN => n51);
   U349 : INV_X1 port map( A => n37, ZN => n85);
   U350 : NAND3_X1 port map( A1 => n35, A2 => n75, A3 => n14, ZN => n45);
   U351 : NAND3_X1 port map( A1 => n44, A2 => n10, A3 => n37, ZN => n116);
   U352 : INV_X1 port map( A => n32, ZN => n52);
   U353 : NAND3_X1 port map( A1 => n124, A2 => n125, A3 => n126, ZN => n89);
   U354 : NAND3_X1 port map( A1 => n136, A2 => n34, A3 => n87, ZN => n133);
   U355 : INV_X1 port map( A => n137, ZN => n136);
   U356 : NAND3_X1 port map( A1 => n66, A2 => n61, A3 => n144, ZN => n122);
   U357 : INV_X1 port map( A => n145, ZN => n144);
   U358 : NAND3_X1 port map( A1 => n151, A2 => n159, A3 => n392, ZN => n156);
   U359 : NAND3_X1 port map( A1 => n147, A2 => n146, A3 => n152, ZN => n155);
   U360 : NAND3_X1 port map( A1 => n174, A2 => n175, A3 => n176, ZN => n173);
   U361 : NAND2_X2 port map( A1 => n177, A2 => n178, ZN => n37);
   U362 : NAND3_X1 port map( A1 => n147, A2 => n179, A3 => n180, ZN => n175);
   U363 : NAND3_X1 port map( A1 => n180, A2 => n147, A3 => n182, ZN => n174);
   U364 : NAND3_X1 port map( A1 => n184, A2 => n185, A3 => n186, ZN => n183);
   U365 : INV_X1 port map( A => n151, ZN => n187);
   U366 : NAND3_X1 port map( A1 => n194, A2 => n195, A3 => n147, ZN => n170);
   U367 : NAND3_X1 port map( A1 => n200, A2 => n146, A3 => n201, ZN => n196);
   U368 : NOR2_X1 port map( A1 => n214, A2 => n215, ZN => GE);
   U369 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n219, ZN
                           => n215);
   U370 : NAND2_X1 port map( A1 => n220, A2 => n221, ZN => n219);
   U371 : NAND3_X1 port map( A1 => n225, A2 => n226, A3 => n227, ZN => n223);
   U372 : NAND2_X1 port map( A1 => n240, A2 => n75, ZN => n235);
   U373 : NAND2_X1 port map( A1 => n242, A2 => n12, ZN => n240);
   U374 : NAND3_X1 port map( A1 => n245, A2 => n48, A3 => n14, ZN => n233);
   U375 : NOR2_X1 port map( A1 => n243, A2 => n249, ZN => n248);
   U376 : INV_X1 port map( A => n112, ZN => n243);
   U377 : NAND3_X1 port map( A1 => n145, A2 => n253, A3 => n254, ZN => n252);
   U378 : NAND2_X1 port map( A1 => n258, A2 => n73, ZN => n257);
   U379 : INV_X1 port map( A => n259, ZN => n258);
   U380 : NAND3_X1 port map( A1 => n121, A2 => n14, A3 => n12, ZN => n260);
   U381 : NAND2_X1 port map( A1 => n261, A2 => n262, ZN => n217);
   U382 : NAND3_X1 port map( A1 => n121, A2 => n14, A3 => n12, ZN => n263);
   U383 : NAND2_X1 port map( A1 => n269, A2 => n270, ZN => n216);
   U384 : NAND2_X1 port map( A1 => n13, A2 => n121, ZN => n271);
   U385 : NAND3_X1 port map( A1 => n274, A2 => n226, A3 => n275, ZN => n272);
   U386 : OAI211_X1 port map( C1 => n276, C2 => n277, A => n278, B => n279, ZN 
                           => n214);
   U387 : INV_X1 port map( A => n286, ZN => n285);
   U388 : NAND2_X1 port map( A1 => n13, A2 => n121, ZN => n287);
   U389 : NAND2_X1 port map( A1 => n290, A2 => n291, ZN => n289);
   U390 : INV_X1 port map( A => n224, ZN => n291);
   U391 : INV_X1 port map( A => n292, ZN => n290);
   U392 : NAND3_X1 port map( A1 => n121, A2 => n14, A3 => n13, ZN => n298);
   U393 : NAND2_X1 port map( A1 => n299, A2 => n300, ZN => n297);
   U394 : NAND3_X1 port map( A1 => n135, A2 => n118, A3 => n64, ZN => n303);
   U395 : INV_X1 port map( A => n87, ZN => n267);
   U396 : NAND3_X1 port map( A1 => n121, A2 => n14, A3 => n119, ZN => n306);
   U397 : NAND2_X1 port map( A1 => n308, A2 => n309, ZN => n305);
   U398 : NAND3_X1 port map( A1 => n135, A2 => n118, A3 => n72, ZN => n312);
   U399 : INV_X1 port map( A => n67, ZN => n134);
   U400 : INV_X1 port map( A => n105, ZN => n118);
   U401 : INV_X1 port map( A => n229, ZN => n135);
   U402 : NAND3_X1 port map( A1 => n315, A2 => n316, A3 => n317, ZN => n277);
   U403 : NAND2_X1 port map( A1 => n325, A2 => n8, ZN => n320);
   U404 : INV_X1 port map( A => n307, ZN => n331);
   U405 : NOR2_X1 port map( A1 => n337, A2 => n6, ZN => n334);
   U406 : INV_X1 port map( A => n244, ZN => n344);
   U407 : INV_X1 port map( A => n114, ZN => n349);
   U408 : NAND3_X1 port map( A1 => n140, A2 => n273, A3 => n3, ZN => n354);
   U409 : INV_X1 port map( A => n48, ZN => n249);
   U410 : NAND2_X1 port map( A1 => n364, A2 => n254, ZN => n362);
   U411 : INV_X1 port map( A => n62, ZN => n364);
   U412 : NAND3_X1 port map( A1 => n368, A2 => n366, A3 => n367, ZN => n276);
   U413 : AOI21_X1 port map( B1 => n369, B2 => n370, A => n371, ZN => n368);
   U414 : NAND3_X1 port map( A1 => n123, A2 => n180, A3 => n87, ZN => n371);
   U415 : NAND3_X1 port map( A1 => n199, A2 => n211, A3 => n200, ZN => n376);
   U416 : NOR2_X1 port map( A1 => n381, A2 => n382, ZN => n369);
   U417 : NAND4_X1 port map( A1 => n383, A2 => n384, A3 => n385, A4 => n386, ZN
                           => n382);
   U418 : NOR2_X1 port map( A1 => n198, A2 => n387, ZN => n385);
   U419 : INV_X1 port map( A => n171, ZN => n387);
   U420 : INV_X1 port map( A => n206, ZN => n198);
   U421 : NAND2_X1 port map( A1 => n390, A2 => n200, ZN => n384);
   U422 : INV_X1 port map( A => n207, ZN => n390);
   U423 : NOR2_X1 port map( A1 => n392, A2 => n327, ZN => n383);
   U424 : NAND3_X1 port map( A1 => n402, A2 => n403, A3 => n404, ZN => n401);
   U425 : NOR2_X1 port map( A1 => n337, A2 => n327, ZN => n404);
   U426 : NOR2_X1 port map( A1 => n405, A2 => n392, ZN => n403);
   U427 : INV_X1 port map( A => n160, ZN => n392);
   U428 : INV_X1 port map( A => n386, ZN => n405);
   U429 : NAND3_X1 port map( A1 => n213, A2 => n417, A3 => n418, ZN => n416);
   U430 : INV_X1 port map( A => n193, ZN => n418);
   U431 : INV_X1 port map( A => n106, ZN => n44);
   U432 : NOR2_X1 port map( A1 => n426, A2 => n361, ZN => n424);
   U433 : INV_X1 port map( A => n36, ZN => n361);
   U434 : INV_X1 port map( A => n254, ZN => n426);
   U435 : NAND3_X1 port map( A1 => n158, A2 => n148, A3 => n430, ZN => n429);
   U436 : NOR2_X1 port map( A1 => n337, A2 => n327, ZN => n430);
   U437 : INV_X1 port map( A => n323, ZN => n327);
   U438 : INV_X1 port map( A => n394, ZN => n337);
   U439 : NAND3_X1 port map( A1 => n417, A2 => n181, A3 => n213, ZN => n326);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_add_2 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end ALU_N32_DW01_add_2;

architecture SYN_cla of ALU_N32_DW01_add_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n39, A2 => n264, ZN => n1);
   U3 : AOI21_X1 port map( B1 => n254, B2 => n253, A => n255, ZN => n2);
   U4 : NOR2_X1 port map( A1 => n16, A2 => n248, ZN => n236);
   U5 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => n55);
   U6 : AND2_X1 port map( A1 => n63, A2 => n56, ZN => n3);
   U7 : AND2_X1 port map( A1 => n188, A2 => n189, ZN => n4);
   U8 : AND2_X1 port map( A1 => n245, A2 => n246, ZN => n5);
   U9 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n72);
   U10 : OAI21_X1 port map( B1 => n265, B2 => n251, A => n252, ZN => n6);
   U11 : INV_X1 port map( A => n6, ZN => n32);
   U12 : AOI21_X1 port map( B1 => n236, B2 => n237, A => n238, ZN => n7);
   U13 : AND2_X2 port map( A1 => n234, A2 => n23, ZN => n8);
   U14 : CLKBUF_X1 port map( A => A(8), Z => n9);
   U15 : AND4_X1 port map( A1 => n85, A2 => n79, A3 => n69, A4 => n72, ZN => 
                           n10);
   U16 : CLKBUF_X1 port map( A => n296, Z => n11);
   U17 : CLKBUF_X1 port map( A => n8, Z => n12);
   U18 : CLKBUF_X1 port map( A => n35, Z => n13);
   U19 : OAI21_X1 port map( B1 => n8, B2 => n226, A => n227, ZN => n14);
   U20 : AOI21_X1 port map( B1 => n236, B2 => n237, A => n238, ZN => n23);
   U21 : NAND2_X1 port map( A1 => n54, A2 => n310, ZN => n15);
   U22 : CLKBUF_X1 port map( A => n239, Z => n16);
   U23 : NAND2_X1 port map( A1 => n306, A2 => n62, ZN => n305);
   U24 : NAND2_X1 port map( A1 => n175, A2 => n176, ZN => n17);
   U25 : AND2_X1 port map( A1 => n32, A2 => n23, ZN => n18);
   U26 : AND3_X1 port map( A1 => n19, A2 => n20, A3 => n89, ZN => n307);
   U27 : NAND3_X1 port map( A1 => n15, A2 => n271, A3 => n308, ZN => n19);
   U28 : AND2_X1 port map( A1 => n88, A2 => n37, ZN => n20);
   U29 : OAI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n21);
   U30 : OAI211_X1 port map( C1 => n12, C2 => n107, A => n111, B => n110, ZN =>
                           n22);
   U31 : AOI21_X1 port map( B1 => n236, B2 => n237, A => n238, ZN => n235);
   U32 : CLKBUF_X1 port map( A => n74, Z => n24);
   U33 : OR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n25);
   U34 : OR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n243);
   U35 : INV_X1 port map( A => A(2), ZN => n26);
   U36 : BUF_X1 port map( A => B(2), Z => n27);
   U37 : NAND2_X1 port map( A1 => n57, A2 => n3, ZN => n302);
   U38 : AND2_X1 port map( A1 => n59, A2 => n296, ZN => n295);
   U39 : OR2_X2 port map( A1 => B(15), A2 => A(15), ZN => n263);
   U40 : OR2_X2 port map( A1 => A(8), A2 => B(8), ZN => n59);
   U41 : NAND2_X1 port map( A1 => n298, A2 => n25, ZN => n300);
   U42 : NAND2_X1 port map( A1 => n299, A2 => n11, ZN => n304);
   U43 : BUF_X1 port map( A => B(0), Z => n28);
   U44 : BUF_X1 port map( A => n261, Z => n29);
   U45 : NOR2_X1 port map( A1 => B(14), A2 => A(14), ZN => n30);
   U46 : AND2_X1 port map( A1 => n243, A2 => n31, ZN => n294);
   U47 : OR2_X1 port map( A1 => A(9), A2 => B(9), ZN => n31);
   U48 : NOR2_X1 port map( A1 => n249, A2 => n250, ZN => n234);
   U49 : OAI21_X1 port map( B1 => n48, B2 => n87, A => n88, ZN => n33);
   U50 : OAI21_X1 port map( B1 => n48, B2 => n87, A => n88, ZN => n84);
   U51 : NAND2_X1 port map( A1 => n32, A2 => n235, ZN => n34);
   U52 : NAND2_X1 port map( A1 => n32, A2 => n7, ZN => n35);
   U53 : NAND2_X1 port map( A1 => n234, A2 => n7, ZN => n108);
   U54 : INV_X1 port map( A => B(2), ZN => n36);
   U55 : NAND2_X1 port map( A1 => n27, A2 => A(2), ZN => n37);
   U56 : INV_X1 port map( A => n34, ZN => n38);
   U57 : AND2_X1 port map( A1 => n295, A2 => n294, ZN => n39);
   U58 : XNOR2_X1 port map( A => n304, B => n40, ZN => SUM(10));
   U59 : NAND2_X1 port map( A1 => n63, A2 => n305, ZN => n40);
   U60 : XNOR2_X1 port map( A => n55, B => n41, ZN => SUM(9));
   U61 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => n41);
   U62 : XOR2_X1 port map( A => n42, B => n278, Z => SUM(13));
   U63 : AND2_X1 port map( A1 => n29, A2 => n260, ZN => n42);
   U64 : AND2_X1 port map( A1 => n219, A2 => n311, ZN => SUM(0));
   U65 : XNOR2_X1 port map( A => n44, B => n300, ZN => SUM(11));
   U66 : NAND2_X1 port map( A1 => n301, A2 => n299, ZN => n44);
   U67 : NOR2_X1 port map( A1 => n38, A2 => n107, ZN => n106);
   U68 : OR2_X2 port map( A1 => n307, A2 => n45, ZN => n61);
   U69 : OR2_X1 port map( A1 => n87, A2 => n273, ZN => n45);
   U70 : AND2_X1 port map( A1 => n146, A2 => n160, ZN => n175);
   U71 : INV_X1 port map( A => n159, ZN => n177);
   U72 : OAI21_X1 port map( B1 => n133, B2 => n130, A => n126, ZN => n132);
   U73 : AND2_X1 port map( A1 => n149, A2 => n47, ZN => n46);
   U74 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => n96);
   U75 : NAND2_X1 port map( A1 => n15, A2 => n121, ZN => n118);
   U76 : NAND2_X1 port map( A1 => n149, A2 => n47, ZN => n159);
   U77 : NAND2_X1 port map( A1 => n46, A2 => n51, ZN => n107);
   U78 : NAND2_X1 port map( A1 => n15, A2 => n119, ZN => n218);
   U79 : NAND2_X1 port map( A1 => n178, A2 => n47, ZN => n160);
   U80 : NAND2_X1 port map( A1 => n51, A2 => n128, ZN => n111);
   U81 : NAND2_X1 port map( A1 => n155, A2 => n156, ZN => n154);
   U82 : NAND2_X1 port map( A1 => n283, A2 => n284, ZN => n278);
   U83 : NAND2_X1 port map( A1 => n285, A2 => n286, ZN => n283);
   U84 : NAND2_X1 port map( A1 => n282, A2 => n267, ZN => n276);
   U85 : AOI21_X1 port map( B1 => n228, B2 => n210, A => n229, ZN => n227);
   U86 : NAND2_X1 port map( A1 => n210, A2 => n217, ZN => n226);
   U87 : AND4_X1 port map( A1 => n179, A2 => n180, A3 => n181, A4 => n182, ZN 
                           => n47);
   U88 : OAI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n70);
   U89 : AND2_X1 port map( A1 => n247, A2 => n72, ZN => n237);
   U90 : OAI21_X1 port map( B1 => n297, B2 => n242, A => n25, ZN => n287);
   U91 : AOI21_X1 port map( B1 => n63, B2 => n56, A => n244, ZN => n297);
   U92 : NAND4_X1 port map( A1 => n217, A2 => n210, A3 => n211, A4 => n147, ZN 
                           => n195);
   U93 : NAND2_X1 port map( A1 => n181, A2 => n187, ZN => n197);
   U94 : XNOR2_X1 port map( A => n169, B => n170, ZN => SUM(25));
   U95 : NOR2_X1 port map( A1 => n171, A2 => n172, ZN => n170);
   U96 : AOI21_X1 port map( B1 => n17, B2 => n144, A => n173, ZN => n169);
   U97 : OAI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n126);
   U98 : NAND2_X1 port map( A1 => n137, A2 => n138, ZN => n135);
   U99 : NOR2_X1 port map( A1 => n49, A2 => n139, ZN => n134);
   U100 : NAND2_X1 port map( A1 => n140, A2 => n141, ZN => n139);
   U101 : AND3_X1 port map( A1 => n90, A2 => n89, A3 => n37, ZN => n48);
   U102 : NAND4_X1 port map( A1 => n266, A2 => n267, A3 => n261, A4 => n263, ZN
                           => n239);
   U103 : NAND4_X1 port map( A1 => n144, A2 => n140, A3 => n141, A4 => n136, ZN
                           => n130);
   U104 : NAND4_X1 port map( A1 => n85, A2 => n79, A3 => n69, A4 => n72, ZN => 
                           n273);
   U105 : NAND2_X1 port map( A1 => n217, A2 => n214, ZN => n233);
   U106 : NAND2_X1 port map( A1 => n144, A2 => n143, ZN => n174);
   U107 : NAND2_X1 port map( A1 => n211, A2 => n216, ZN => n225);
   U108 : NAND2_X1 port map( A1 => n210, A2 => n213, ZN => n230);
   U109 : NAND2_X1 port map( A1 => n180, A2 => n188, ZN => n202);
   U110 : NAND2_X1 port map( A1 => n179, A2 => n189, ZN => n206);
   U111 : NAND2_X1 port map( A1 => n319, A2 => n67, ZN => n73);
   U112 : NAND2_X1 port map( A1 => n136, A2 => n137, ZN => n151);
   U113 : OAI21_X1 port map( B1 => n152, B2 => n153, A => n138, ZN => n150);
   U114 : NAND2_X1 port map( A1 => n154, A2 => n141, ZN => n153);
   U115 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => n65);
   U116 : NAND2_X1 port map( A1 => n68, A2 => n67, ZN => n66);
   U117 : NAND2_X1 port map( A1 => n70, A2 => n69, ZN => n68);
   U118 : NOR2_X1 port map( A1 => n163, A2 => n164, ZN => n162);
   U119 : NAND2_X1 port map( A1 => n312, A2 => n313, ZN => n69);
   U120 : NAND2_X1 port map( A1 => n72, A2 => n247, ZN => n60);
   U121 : NAND2_X1 port map( A1 => n298, A2 => n299, ZN => n242);
   U122 : OAI21_X1 port map( B1 => n100, B2 => n101, A => n102, ZN => n98);
   U123 : NAND2_X1 port map( A1 => n103, A2 => n104, ZN => n101);
   U124 : NOR2_X1 port map( A1 => n106, A2 => n105, ZN => n100);
   U125 : XNOR2_X1 port map( A => n64, B => n58, ZN => SUM(8));
   U126 : XNOR2_X1 port map( A => n190, B => n191, ZN => SUM(23));
   U127 : NAND2_X1 port map( A1 => n182, A2 => n186, ZN => n191);
   U128 : OAI21_X1 port map( B1 => n193, B2 => n50, A => n194, ZN => n192);
   U129 : XNOR2_X1 port map( A => n279, B => n280, ZN => SUM(14));
   U130 : NOR2_X1 port map( A1 => n281, A2 => n30, ZN => n280);
   U131 : AOI21_X1 port map( B1 => n29, B2 => n278, A => n282, ZN => n279);
   U132 : XNOR2_X1 port map( A => n289, B => n290, ZN => SUM(12));
   U133 : NOR2_X1 port map( A1 => n288, A2 => n291, ZN => n290);
   U134 : NOR2_X1 port map( A1 => n292, A2 => n293, ZN => n289);
   U135 : OAI21_X1 port map( B1 => n241, B2 => n242, A => n25, ZN => n240);
   U136 : NOR2_X1 port map( A1 => n5, A2 => n244, ZN => n241);
   U137 : NAND2_X1 port map( A1 => n57, A2 => n56, ZN => n306);
   U138 : NAND2_X1 port map( A1 => n168, A2 => n140, ZN => n156);
   U139 : NAND2_X1 port map( A1 => n142, A2 => n143, ZN => n168);
   U140 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => n146);
   U141 : OAI21_X1 port map( B1 => n4, B2 => n184, A => n185, ZN => n183);
   U142 : AND2_X1 port map( A1 => n186, A2 => n187, ZN => n185);
   U143 : NOR2_X1 port map( A1 => n78, A2 => n75, ZN => n77);
   U144 : INV_X1 port map( A => n219, ZN => n121);
   U145 : NAND2_X1 port map( A1 => n125, A2 => n127, ZN => n131);
   U146 : NAND2_X1 port map( A1 => n54, A2 => n310, ZN => n120);
   U147 : AND2_X1 port map( A1 => n142, A2 => n143, ZN => n49);
   U148 : NAND2_X1 port map( A1 => n144, A2 => n140, ZN => n155);
   U149 : NAND2_X1 port map( A1 => n71, A2 => n67, ZN => n321);
   U150 : NAND2_X1 port map( A1 => n314, A2 => n315, ZN => n79);
   U151 : NAND2_X1 port map( A1 => n145, A2 => n146, ZN => n128);
   U152 : NAND2_X1 port map( A1 => n104, A2 => n109, ZN => n123);
   U153 : NAND2_X1 port map( A1 => n208, A2 => n209, ZN => n148);
   U154 : AND2_X1 port map( A1 => n215, A2 => n216, ZN => n208);
   U155 : NAND2_X1 port map( A1 => n213, A2 => n214, ZN => n212);
   U156 : NAND2_X1 port map( A1 => n97, A2 => n88, ZN => n92);
   U157 : NAND2_X1 port map( A1 => n147, A2 => n215, ZN => n220);
   U158 : AND3_X1 port map( A1 => n34, A2 => n149, A3 => n179, ZN => n50);
   U159 : NAND2_X1 port map( A1 => n256, A2 => n263, ZN => n274);
   U160 : NAND2_X1 port map( A1 => n178, A2 => n179, ZN => n196);
   U161 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => n112);
   U162 : NAND2_X1 port map( A1 => n148, A2 => n147, ZN => n205);
   U163 : NAND2_X1 port map( A1 => n124, A2 => n125, ZN => n110);
   U164 : NAND2_X1 port map( A1 => n52, A2 => n325, ZN => n311);
   U165 : NAND2_X1 port map( A1 => n180, A2 => n181, ZN => n184);
   U166 : NAND2_X1 port map( A1 => n83, A2 => n85, ZN => n86);
   U167 : NAND2_X1 port map( A1 => n314, A2 => n315, ZN => n318);
   U168 : NAND2_X1 port map( A1 => n312, A2 => n313, ZN => n319);
   U169 : AND2_X1 port map( A1 => n129, A2 => n125, ZN => n51);
   U170 : AND2_X1 port map( A1 => n180, A2 => n181, ZN => n194);
   U171 : AND2_X1 port map( A1 => n189, A2 => n196, ZN => n203);
   U172 : AND2_X1 port map( A1 => n11, A2 => n62, ZN => n303);
   U173 : INV_X1 port map( A => n2, ZN => n250);
   U174 : AOI21_X1 port map( B1 => n254, B2 => n253, A => n255, ZN => n252);
   U175 : XNOR2_X1 port map( A => n131, B => n132, ZN => SUM(28));
   U176 : XNOR2_X1 port map( A => n117, B => n96, ZN => SUM(2));
   U177 : NAND2_X1 port map( A1 => B(24), A2 => A(24), ZN => n143);
   U178 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n99);
   U179 : OR2_X1 port map( A1 => B(17), A2 => A(17), ZN => n210);
   U180 : OR2_X1 port map( A1 => A(10), A2 => B(10), ZN => n296);
   U181 : OR2_X1 port map( A1 => B(13), A2 => A(13), ZN => n261);
   U182 : OR2_X1 port map( A1 => B(20), A2 => A(20), ZN => n179);
   U183 : NAND2_X1 port map( A1 => B(23), A2 => A(23), ZN => n186);
   U184 : OAI211_X1 port map( C1 => n257, C2 => n258, A => n259, B => n260, ZN 
                           => n254);
   U185 : OR2_X1 port map( A1 => B(19), A2 => A(19), ZN => n147);
   U186 : OR2_X1 port map( A1 => B(22), A2 => A(22), ZN => n181);
   U187 : OR2_X1 port map( A1 => B(24), A2 => A(24), ZN => n144);
   U188 : OR2_X1 port map( A1 => B(28), A2 => A(28), ZN => n125);
   U189 : OR2_X1 port map( A1 => B(16), A2 => A(16), ZN => n217);
   U190 : OR2_X1 port map( A1 => B(26), A2 => A(26), ZN => n141);
   U191 : OR2_X1 port map( A1 => B(23), A2 => A(23), ZN => n182);
   U192 : OR2_X1 port map( A1 => B(27), A2 => A(27), ZN => n136);
   U193 : OR2_X1 port map( A1 => B(18), A2 => A(18), ZN => n211);
   U194 : OR2_X1 port map( A1 => B(29), A2 => A(29), ZN => n104);
   U195 : XNOR2_X1 port map( A => n218, B => n121, ZN => SUM(1));
   U196 : OR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n62);
   U197 : NOR2_X1 port map( A1 => n323, A2 => n324, ZN => n322);
   U198 : OR2_X1 port map( A1 => B(4), A2 => A(4), ZN => n85);
   U199 : OR2_X1 port map( A1 => B(21), A2 => A(21), ZN => n180);
   U200 : OR2_X1 port map( A1 => A(14), A2 => B(14), ZN => n267);
   U201 : OR2_X1 port map( A1 => B(25), A2 => A(25), ZN => n140);
   U202 : OR2_X1 port map( A1 => B(3), A2 => A(3), ZN => n97);
   U203 : OR2_X1 port map( A1 => B(30), A2 => A(30), ZN => n103);
   U204 : NAND2_X1 port map( A1 => n316, A2 => n317, ZN => n247);
   U205 : NOR2_X1 port map( A1 => n321, A2 => n322, ZN => n316);
   U206 : OR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n266);
   U207 : NOR2_X1 port map( A1 => n157, A2 => n158, ZN => n152);
   U208 : NAND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n83);
   U209 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n320);
   U210 : NAND2_X1 port map( A1 => B(28), A2 => A(28), ZN => n127);
   U211 : NAND2_X1 port map( A1 => B(29), A2 => A(29), ZN => n109);
   U212 : NAND2_X1 port map( A1 => B(17), A2 => A(17), ZN => n213);
   U213 : NAND2_X1 port map( A1 => B(16), A2 => A(16), ZN => n214);
   U214 : NAND2_X1 port map( A1 => B(21), A2 => A(21), ZN => n188);
   U215 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => n57);
   U216 : NAND2_X1 port map( A1 => n56, A2 => n59, ZN => n64);
   U217 : NAND2_X1 port map( A1 => B(30), A2 => A(30), ZN => n102);
   U218 : NAND2_X1 port map( A1 => B(20), A2 => A(20), ZN => n189);
   U219 : NAND2_X1 port map( A1 => B(27), A2 => A(27), ZN => n137);
   U220 : NAND2_X1 port map( A1 => B(26), A2 => A(26), ZN => n138);
   U221 : INV_X1 port map( A => B(5), ZN => n314);
   U222 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n63);
   U223 : OAI211_X1 port map( C1 => A(2), C2 => n27, A => A(1), B => n53, ZN =>
                           n89);
   U224 : INV_X1 port map( A => A(2), ZN => n309);
   U225 : NAND2_X1 port map( A1 => B(19), A2 => A(19), ZN => n215);
   U226 : NAND2_X1 port map( A1 => B(25), A2 => A(25), ZN => n142);
   U227 : OAI22_X1 port map( A1 => A(10), A2 => B(10), B1 => A(9), B2 => B(9), 
                           ZN => n244);
   U228 : NAND2_X1 port map( A1 => A(10), A2 => B(10), ZN => n299);
   U229 : NAND2_X1 port map( A1 => B(18), A2 => A(18), ZN => n216);
   U230 : NAND2_X1 port map( A1 => B(13), A2 => A(13), ZN => n260);
   U231 : NAND2_X1 port map( A1 => B(15), A2 => A(15), ZN => n256);
   U232 : INV_X1 port map( A => B(6), ZN => n312);
   U233 : XNOR2_X1 port map( A => n66, B => n65, ZN => SUM(7));
   U234 : OAI21_X1 port map( B1 => n226, B2 => n8, A => n227, ZN => n224);
   U235 : OAI211_X1 port map( C1 => n8, C2 => n107, A => n111, B => n110, ZN =>
                           n116);
   U236 : XNOR2_X1 port map( A => n13, B => n233, ZN => SUM(16));
   U237 : AOI21_X1 port map( B1 => n35, B2 => n46, A => n128, ZN => n133);
   U238 : NAND2_X1 port map( A1 => n35, A2 => n177, ZN => n176);
   U239 : NAND2_X1 port map( A1 => B(22), A2 => A(22), ZN => n187);
   U240 : NAND2_X1 port map( A1 => n203, A2 => n204, ZN => n201);
   U241 : AOI21_X1 port map( B1 => n248, B2 => n287, A => n288, ZN => n285);
   U242 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n71);
   U243 : NAND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n284);
   U244 : NOR2_X1 port map( A1 => n265, A2 => n1, ZN => n249);
   U245 : XNOR2_X1 port map( A => n274, B => n275, ZN => SUM(15));
   U246 : NOR2_X1 port map( A1 => n18, A2 => n159, ZN => n158);
   U247 : XNOR2_X1 port map( A => n150, B => n151, ZN => SUM(27));
   U248 : XNOR2_X1 port map( A => n98, B => n99, ZN => SUM(31));
   U249 : INV_X1 port map( A => A(5), ZN => n315);
   U250 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => n76);
   U251 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => n88);
   U252 : NAND2_X1 port map( A1 => n192, A2 => n187, ZN => n190);
   U253 : NAND2_X1 port map( A1 => n309, A2 => n36, ZN => n122);
   U254 : NAND2_X1 port map( A1 => n36, A2 => n26, ZN => n271);
   U255 : NAND2_X1 port map( A1 => n39, A2 => n264, ZN => n251);
   U256 : NOR2_X1 port map( A1 => n240, A2 => n239, ZN => n238);
   U257 : NAND2_X1 port map( A1 => B(14), A2 => A(14), ZN => n259);
   U258 : NAND2_X1 port map( A1 => n27, A2 => A(2), ZN => n91);
   U259 : AND2_X1 port map( A1 => n88, A2 => n91, ZN => n269);
   U260 : NAND2_X1 port map( A1 => n271, A2 => n37, ZN => n117);
   U261 : INV_X1 port map( A => A(0), ZN => n325);
   U262 : NAND2_X1 port map( A1 => n28, A2 => A(0), ZN => n219);
   U263 : AND2_X1 port map( A1 => n28, A2 => A(0), ZN => n308);
   U264 : AND2_X1 port map( A1 => n28, A2 => A(0), ZN => n272);
   U265 : NAND2_X1 port map( A1 => B(8), A2 => n9, ZN => n56);
   U266 : OAI21_X1 port map( B1 => n81, B2 => n82, A => n83, ZN => n80);
   U267 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n298);
   U268 : NAND2_X1 port map( A1 => n294, A2 => n295, ZN => n248);
   U269 : AOI21_X1 port map( B1 => n60, B2 => n61, A => n248, ZN => n293);
   U270 : NAND2_X1 port map( A1 => n302, A2 => n303, ZN => n301);
   U271 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => n58);
   U272 : AOI21_X1 port map( B1 => n165, B2 => n166, A => n167, ZN => n161);
   U273 : NAND2_X1 port map( A1 => n175, A2 => n176, ZN => n166);
   U274 : NOR2_X1 port map( A1 => A(6), A2 => B(6), ZN => n323);
   U275 : INV_X1 port map( A => A(6), ZN => n313);
   U276 : NAND2_X1 port map( A1 => B(6), A2 => A(6), ZN => n67);
   U277 : XNOR2_X1 port map( A => n161, B => n162, ZN => SUM(26));
   U278 : INV_X1 port map( A => B(1), ZN => n54);
   U279 : NAND2_X1 port map( A1 => n53, A2 => A(1), ZN => n119);
   U280 : INV_X1 port map( A => A(1), ZN => n310);
   U281 : INV_X1 port map( A => B(0), ZN => n52);
   U282 : INV_X1 port map( A => n54, ZN => n53);
   U283 : XNOR2_X1 port map( A => n21, B => n73, ZN => SUM(6));
   U284 : XNOR2_X1 port map( A => n24, B => n77, ZN => SUM(5));
   U285 : INV_X1 port map( A => n79, ZN => n75);
   U286 : INV_X1 port map( A => n76, ZN => n78);
   U287 : INV_X1 port map( A => n80, ZN => n74);
   U288 : INV_X1 port map( A => n84, ZN => n82);
   U289 : INV_X1 port map( A => n85, ZN => n81);
   U290 : XNOR2_X1 port map( A => n86, B => n33, ZN => SUM(4));
   U291 : XNOR2_X1 port map( A => n92, B => n93, ZN => SUM(3));
   U292 : OAI21_X1 port map( B1 => n94, B2 => n95, A => n37, ZN => n93);
   U293 : INV_X1 port map( A => n96, ZN => n94);
   U294 : NAND3_X1 port map( A1 => n109, A2 => n110, A3 => n111, ZN => n105);
   U295 : XNOR2_X1 port map( A => n113, B => n112, ZN => SUM(30));
   U296 : OAI21_X1 port map( B1 => n114, B2 => n115, A => n109, ZN => n113);
   U297 : INV_X1 port map( A => n104, ZN => n115);
   U298 : INV_X1 port map( A => n116, ZN => n114);
   U299 : XNOR2_X1 port map( A => n22, B => n123, ZN => SUM(29));
   U300 : NAND2_X1 port map( A1 => n126, A2 => n127, ZN => n124);
   U301 : INV_X1 port map( A => n130, ZN => n129);
   U302 : NAND3_X1 port map( A1 => n47, A2 => n147, A3 => n148, ZN => n145);
   U303 : NAND3_X1 port map( A1 => n156, A2 => n146, A3 => n160, ZN => n157);
   U304 : INV_X1 port map( A => n141, ZN => n164);
   U305 : INV_X1 port map( A => n138, ZN => n163);
   U306 : INV_X1 port map( A => n156, ZN => n167);
   U307 : INV_X1 port map( A => n155, ZN => n165);
   U308 : INV_X1 port map( A => n140, ZN => n172);
   U309 : INV_X1 port map( A => n142, ZN => n171);
   U310 : INV_X1 port map( A => n143, ZN => n173);
   U311 : XNOR2_X1 port map( A => n17, B => n174, ZN => SUM(24));
   U312 : NAND3_X1 port map( A1 => n188, A2 => n189, A3 => n196, ZN => n193);
   U313 : XNOR2_X1 port map( A => n198, B => n197, ZN => SUM(22));
   U314 : OAI21_X1 port map( B1 => n199, B2 => n200, A => n188, ZN => n198);
   U315 : INV_X1 port map( A => n180, ZN => n200);
   U316 : INV_X1 port map( A => n201, ZN => n199);
   U317 : XNOR2_X1 port map( A => n202, B => n201, ZN => SUM(21));
   U318 : NAND3_X1 port map( A1 => n108, A2 => n149, A3 => n179, ZN => n204);
   U319 : INV_X1 port map( A => n195, ZN => n149);
   U320 : INV_X1 port map( A => n205, ZN => n178);
   U321 : XNOR2_X1 port map( A => n206, B => n207, ZN => SUM(20));
   U322 : OAI21_X1 port map( B1 => n18, B2 => n195, A => n205, ZN => n207);
   U323 : NAND3_X1 port map( A1 => n210, A2 => n211, A3 => n212, ZN => n209);
   U324 : XNOR2_X1 port map( A => n221, B => n220, ZN => SUM(19));
   U325 : OAI21_X1 port map( B1 => n222, B2 => n223, A => n216, ZN => n221);
   U326 : INV_X1 port map( A => n211, ZN => n223);
   U327 : INV_X1 port map( A => n14, ZN => n222);
   U328 : XNOR2_X1 port map( A => n224, B => n225, ZN => SUM(18));
   U329 : INV_X1 port map( A => n213, ZN => n229);
   U330 : INV_X1 port map( A => n214, ZN => n228);
   U331 : XNOR2_X1 port map( A => n230, B => n231, ZN => SUM(17));
   U332 : OAI21_X1 port map( B1 => n18, B2 => n232, A => n214, ZN => n231);
   U333 : INV_X1 port map( A => n217, ZN => n232);
   U334 : NAND2_X1 port map( A1 => A(8), A2 => B(8), ZN => n246);
   U335 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n245);
   U336 : INV_X1 port map( A => n256, ZN => n255);
   U337 : NAND2_X1 port map( A1 => A(12), A2 => B(12), ZN => n258);
   U338 : INV_X1 port map( A => n261, ZN => n257);
   U339 : NOR2_X1 port map( A1 => n262, A2 => n30, ZN => n253);
   U340 : INV_X1 port map( A => n263, ZN => n262);
   U341 : INV_X1 port map( A => n239, ZN => n264);
   U342 : NAND3_X1 port map( A1 => n268, A2 => n97, A3 => n10, ZN => n265);
   U343 : NAND3_X1 port map( A1 => n270, A2 => n269, A3 => n89, ZN => n268);
   U344 : NAND3_X1 port map( A1 => n122, A2 => n120, A3 => n272, ZN => n270);
   U345 : NAND3_X1 port map( A1 => n259, A2 => n276, A3 => n277, ZN => n275);
   U346 : NAND3_X1 port map( A1 => n278, A2 => n267, A3 => n29, ZN => n277);
   U347 : INV_X1 port map( A => n259, ZN => n281);
   U348 : INV_X1 port map( A => n260, ZN => n282);
   U349 : NAND3_X1 port map( A1 => n60, A2 => n287, A3 => n61, ZN => n286);
   U350 : INV_X1 port map( A => n284, ZN => n291);
   U351 : INV_X1 port map( A => n266, ZN => n288);
   U352 : INV_X1 port map( A => n287, ZN => n292);
   U353 : NAND3_X1 port map( A1 => n15, A2 => n122, A3 => n308, ZN => n90);
   U354 : INV_X1 port map( A => n271, ZN => n95);
   U355 : INV_X1 port map( A => n97, ZN => n87);
   U356 : NAND3_X1 port map( A1 => n318, A2 => n319, A3 => n320, ZN => n317);
   U357 : NAND2_X1 port map( A1 => A(5), A2 => B(5), ZN => n324);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_sub_2 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end ALU_N32_DW01_sub_2;

architecture SYN_cla of ALU_N32_DW01_sub_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408 : std_logic;

begin
   
   U3 : AND4_X2 port map( A1 => n271, A2 => n272, A3 => n29, A4 => n269, ZN => 
                           n1);
   U4 : INV_X4 port map( A => n1, ZN => n255);
   U5 : AND2_X2 port map( A1 => B(0), A2 => n394, ZN => n66);
   U6 : AND4_X2 port map( A1 => n356, A2 => n19, A3 => n17, A4 => n81, ZN => 
                           n28);
   U7 : INV_X1 port map( A => n11, ZN => n173);
   U8 : NAND2_X1 port map( A1 => B(21), A2 => n257, ZN => n225);
   U9 : AND2_X1 port map( A1 => n100, A2 => n101, ZN => n44);
   U10 : AND2_X1 port map( A1 => n185, A2 => n205, ZN => n56);
   U11 : AND2_X1 port map( A1 => n32, A2 => n302, ZN => n2);
   U12 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => n118);
   U13 : AND2_X1 port map( A1 => n112, A2 => n113, ZN => n3);
   U14 : AND2_X1 port map( A1 => n294, A2 => B(17), ZN => n4);
   U15 : AND2_X1 port map( A1 => n143, A2 => n5, ZN => n137);
   U16 : AND2_X1 port map( A1 => n141, A2 => n39, ZN => n5);
   U17 : INV_X1 port map( A => n33, ZN => n82);
   U18 : NAND3_X1 port map( A1 => n390, A2 => n16, A3 => n307, ZN => n6);
   U19 : NOR2_X1 port map( A1 => n12, A2 => n13, ZN => n7);
   U20 : CLKBUF_X1 port map( A => n209, Z => n8);
   U21 : NAND2_X1 port map( A1 => B(6), A2 => n399, ZN => n9);
   U22 : NAND2_X1 port map( A1 => n53, A2 => n299, ZN => n10);
   U23 : AND2_X1 port map( A1 => B(25), A2 => n201, ZN => n11);
   U24 : AND2_X1 port map( A1 => n378, A2 => A(9), ZN => n367);
   U25 : NOR2_X1 port map( A1 => n12, A2 => n13, ZN => n308);
   U26 : NAND3_X1 port map( A1 => n324, A2 => n109, A3 => n47, ZN => n12);
   U27 : NAND2_X1 port map( A1 => n28, A2 => n40, ZN => n13);
   U28 : INV_X1 port map( A => n44, ZN => n98);
   U29 : CLKBUF_X1 port map( A => A(1), Z => n31);
   U30 : NOR2_X1 port map( A1 => n148, A2 => n66, ZN => n14);
   U31 : XNOR2_X1 port map( A => n132, B => n15, ZN => DIFF(30));
   U32 : NAND2_X1 port map( A1 => n124, A2 => n130, ZN => n15);
   U33 : CLKBUF_X1 port map( A => n212, Z => n16);
   U34 : NAND2_X1 port map( A1 => B(9), A2 => n368, ZN => n17);
   U35 : CLKBUF_X1 port map( A => n9, Z => n18);
   U36 : NAND2_X1 port map( A1 => B(10), A2 => n407, ZN => n19);
   U37 : CLKBUF_X1 port map( A => A(11), Z => n20);
   U38 : INV_X1 port map( A => n31, ZN => n21);
   U39 : NAND3_X1 port map( A1 => n390, A2 => n16, A3 => n307, ZN => n86);
   U40 : CLKBUF_X1 port map( A => n81, Z => n22);
   U41 : CLKBUF_X1 port map( A => n267, Z => n23);
   U42 : AND2_X1 port map( A1 => n326, A2 => n327, ZN => n24);
   U43 : CLKBUF_X1 port map( A => A(0), Z => n25);
   U44 : BUF_X1 port map( A => n218, Z => n26);
   U45 : OAI211_X1 port map( C1 => n366, C2 => n367, A => n19, B => n17, ZN => 
                           n27);
   U46 : NAND2_X1 port map( A1 => n290, A2 => B(18), ZN => n29);
   U47 : AND2_X1 port map( A1 => B(13), A2 => n350, ZN => n30);
   U48 : OAI21_X1 port map( B1 => n24, B2 => n325, A => n212, ZN => n324);
   U49 : NAND2_X1 port map( A1 => n266, A2 => n4, ZN => n265);
   U50 : OR2_X1 port map( A1 => n74, A2 => A(2), ZN => n382);
   U51 : BUF_X1 port map( A => n322, Z => n32);
   U52 : AND2_X1 port map( A1 => n93, A2 => n344, ZN => n33);
   U53 : NAND2_X1 port map( A1 => n53, A2 => n299, ZN => n52);
   U54 : AND2_X1 port map( A1 => n42, A2 => n299, ZN => n34);
   U55 : AND2_X1 port map( A1 => n42, A2 => n299, ZN => n48);
   U56 : OAI211_X1 port map( C1 => n366, C2 => n367, A => n364, B => n365, ZN 
                           => n35);
   U57 : INV_X1 port map( A => n28, ZN => n36);
   U58 : AND2_X1 port map( A1 => B(12), A2 => n360, ZN => n37);
   U59 : AND3_X1 port map( A1 => n383, A2 => n385, A3 => n382, ZN => n38);
   U60 : NAND2_X1 port map( A1 => n317, A2 => n318, ZN => n39);
   U61 : AND4_X1 port map( A1 => n322, A2 => n323, A3 => n306, A4 => n305, ZN 
                           => n40);
   U62 : INV_X1 port map( A => n49, ZN => n41);
   U63 : NOR2_X1 port map( A1 => n7, A2 => n309, ZN => n42);
   U64 : AND2_X1 port map( A1 => n50, A2 => n43, ZN => n138);
   U65 : AND2_X1 port map( A1 => n139, A2 => n140, ZN => n43);
   U66 : XNOR2_X1 port map( A => n248, B => n45, ZN => DIFF(22));
   U67 : AND2_X1 port map( A1 => n226, A2 => n235, ZN => n45);
   U68 : NAND3_X1 port map( A1 => n115, A2 => n114, A3 => n3, ZN => n111);
   U69 : AND2_X1 port map( A1 => n73, A2 => n387, ZN => n46);
   U70 : AND4_X2 port map( A1 => n102, A2 => n91, A3 => n97, A4 => n93, ZN => 
                           n47);
   U71 : AND2_X1 port map( A1 => B(5), A2 => n315, ZN => n49);
   U72 : CLKBUF_X1 port map( A => n220, Z => n50);
   U73 : XNOR2_X1 port map( A => n192, B => n51, ZN => DIFF(26));
   U74 : AND2_X1 port map( A1 => n166, A2 => n170, ZN => n51);
   U75 : NOR2_X1 port map( A1 => n308, A2 => n309, ZN => n53);
   U76 : NOR2_X1 port map( A1 => n157, A2 => n55, ZN => n59);
   U77 : XNOR2_X1 port map( A => n236, B => n54, ZN => DIFF(23));
   U78 : AND2_X1 port map( A1 => n227, A2 => n231, ZN => n54);
   U79 : XOR2_X1 port map( A => n347, B => n348, Z => DIFF(13));
   U80 : AND2_X1 port map( A1 => n94, A2 => n89, ZN => n60);
   U81 : AND2_X1 port map( A1 => B(28), A2 => n176, ZN => n55);
   U82 : INV_X1 port map( A => n121, ZN => n119);
   U83 : AOI21_X1 port map( B1 => n82, B2 => n363, A => n36, ZN => n362);
   U84 : AOI21_X1 port map( B1 => n82, B2 => n363, A => n338, ZN => n351);
   U85 : INV_X1 port map( A => n117, ZN => n116);
   U86 : OAI21_X1 port map( B1 => n56, B2 => n157, A => n162, ZN => n161);
   U87 : NOR2_X1 port map( A1 => n118, A2 => n129, ZN => n126);
   U88 : NOR2_X1 port map( A1 => n338, A2 => n342, ZN => n341);
   U89 : NAND2_X1 port map( A1 => n59, A2 => n155, ZN => n121);
   U90 : NAND2_X1 port map( A1 => n156, A2 => n59, ZN => n117);
   U91 : NOR2_X1 port map( A1 => n122, A2 => n123, ZN => n113);
   U92 : NOR2_X1 port map( A1 => n126, A2 => n127, ZN => n112);
   U93 : NAND2_X1 port map( A1 => n119, A2 => n120, ZN => n114);
   U94 : NAND2_X1 port map( A1 => n1, A2 => n58, ZN => n191);
   U95 : NOR2_X1 port map( A1 => n37, A2 => n353, ZN => n352);
   U96 : INV_X1 port map( A => n118, ZN => n120);
   U97 : NAND2_X1 port map( A1 => n141, A2 => n142, ZN => n309);
   U98 : OAI21_X1 port map( B1 => n254, B2 => n223, A => n224, ZN => n241);
   U99 : OAI21_X1 port map( B1 => n395, B2 => n396, A => n60, ZN => n344);
   U100 : NAND2_X1 port map( A1 => n215, A2 => n216, ZN => n213);
   U101 : OAI21_X1 port map( B1 => n163, B2 => n164, A => n165, ZN => n153);
   U102 : NAND2_X1 port map( A1 => n166, A2 => n167, ZN => n164);
   U103 : NOR2_X1 port map( A1 => n168, A2 => n169, ZN => n163);
   U104 : NAND2_X1 port map( A1 => n170, A2 => n171, ZN => n169);
   U105 : OAI211_X1 port map( C1 => n232, C2 => n233, A => n234, B => n235, ZN 
                           => n229);
   U106 : INV_X1 port map( A => n225, ZN => n233);
   U107 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => n139);
   U108 : AND2_X1 port map( A1 => n305, A2 => n306, ZN => n300);
   U109 : OAI211_X1 port map( C1 => n30, C2 => n302, A => n303, B => n304, ZN 
                           => n301);
   U110 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n117, ZN => n135);
   U111 : NAND4_X1 port map( A1 => n174, A2 => n173, A3 => n166, A4 => n167, ZN
                           => n157);
   U112 : NAND2_X1 port map( A1 => n271, A2 => n267, ZN => n296);
   U113 : NAND2_X1 port map( A1 => n356, A2 => n320, ZN => n370);
   U114 : XOR2_X1 port map( A => n57, B => n332, Z => DIFF(14));
   U115 : AND2_X1 port map( A1 => n306, A2 => n303, ZN => n57);
   U116 : NAND2_X1 port map( A1 => n91, A2 => n89, ZN => n95);
   U117 : NAND2_X1 port map( A1 => n225, A2 => n234, ZN => n252);
   U118 : NAND2_X1 port map( A1 => n224, A2 => n232, ZN => n258);
   U119 : NAND2_X1 port map( A1 => n266, A2 => n29, ZN => n285);
   U120 : NAND2_X1 port map( A1 => n268, A2 => n287, ZN => n286);
   U121 : NAND2_X1 port map( A1 => n173, A2 => n171, ZN => n197);
   U122 : OAI21_X1 port map( B1 => n56, B2 => n199, A => n172, ZN => n198);
   U123 : XOR2_X1 port map( A => n56, B => n202, Z => DIFF(24));
   U124 : NAND2_X1 port map( A1 => n174, A2 => n172, ZN => n202);
   U125 : AOI21_X1 port map( B1 => n339, B2 => n340, A => n341, ZN => n335);
   U126 : OAI21_X1 port map( B1 => n283, B2 => n268, A => n266, ZN => n282);
   U127 : AND4_X1 port map( A1 => n224, A2 => n225, A3 => n226, A4 => n227, ZN 
                           => n58);
   U128 : AOI21_X1 port map( B1 => n212, B2 => n213, A => n214, ZN => n208);
   U129 : NOR2_X1 port map( A1 => n118, A2 => n125, ZN => n122);
   U130 : NOR2_X1 port map( A1 => n11, A2 => n172, ZN => n168);
   U131 : NOR2_X1 port map( A1 => n118, A2 => n128, ZN => n127);
   U132 : NAND2_X1 port map( A1 => n1, A2 => n224, ZN => n247);
   U133 : NOR2_X1 port map( A1 => n351, A2 => n352, ZN => n347);
   U134 : NAND2_X1 port map( A1 => n323, A2 => n304, ZN => n348);
   U135 : OAI21_X1 port map( B1 => n330, B2 => n331, A => n303, ZN => n329);
   U136 : OAI21_X1 port map( B1 => n133, B2 => n134, A => n128, ZN => n132);
   U137 : NOR2_X1 port map( A1 => n135, A2 => n136, ZN => n133);
   U138 : NAND2_X1 port map( A1 => n63, A2 => n121, ZN => n136);
   U139 : AND2_X1 port map( A1 => n174, A2 => n173, ZN => n61);
   U140 : NAND2_X1 port map( A1 => n317, A2 => n318, ZN => n142);
   U141 : NAND2_X1 port map( A1 => n153, A2 => n154, ZN => n129);
   U142 : NAND2_X1 port map( A1 => n209, A2 => n310, ZN => n141);
   U143 : AOI21_X1 port map( B1 => n60, B2 => n311, A => n312, ZN => n310);
   U144 : XNOR2_X1 port map( A => n83, B => n84, ZN => DIFF(8));
   U145 : XNOR2_X1 port map( A => n177, B => n178, ZN => DIFF(27));
   U146 : XOR2_X1 port map( A => n62, B => n374, Z => DIFF(10));
   U147 : AND2_X1 port map( A1 => n364, A2 => n319, ZN => n62);
   U148 : XNOR2_X1 port map( A => n291, B => n292, ZN => DIFF(17));
   U149 : NAND2_X1 port map( A1 => n272, A2 => n268, ZN => n292);
   U150 : NAND2_X1 port map( A1 => n23, A2 => n295, ZN => n291);
   U151 : XNOR2_X1 port map( A => n75, B => n76, ZN => DIFF(9));
   U152 : AOI21_X1 port map( B1 => n80, B2 => n22, A => n68, ZN => n75);
   U153 : XNOR2_X1 port map( A => n358, B => n2, ZN => DIFF(12));
   U154 : NOR2_X1 port map( A1 => n361, A2 => n362, ZN => n358);
   U155 : OAI21_X1 port map( B1 => n241, B2 => n242, A => n243, ZN => n240);
   U156 : NAND2_X1 port map( A1 => n225, A2 => n226, ZN => n242);
   U157 : AOI21_X1 port map( B1 => n244, B2 => n226, A => n245, ZN => n243);
   U158 : OAI21_X1 port map( B1 => n185, B2 => n186, A => n187, ZN => n184);
   U159 : AOI21_X1 port map( B1 => n188, B2 => n166, A => n189, ZN => n187);
   U160 : AND2_X1 port map( A1 => n129, A2 => n125, ZN => n63);
   U161 : NAND2_X1 port map( A1 => n66, A2 => n276, ZN => n150);
   U162 : NAND2_X1 port map( A1 => n377, A2 => n79, ZN => n374);
   U163 : NAND2_X1 port map( A1 => n379, A2 => n380, ZN => n377);
   U164 : NAND2_X1 port map( A1 => n354, A2 => n302, ZN => n340);
   U165 : NAND2_X1 port map( A1 => n355, A2 => n356, ZN => n354);
   U166 : NAND2_X1 port map( A1 => n154, A2 => n125, ZN => n160);
   U167 : NAND2_X1 port map( A1 => n131, A2 => n128, ZN => n151);
   U168 : AND2_X1 port map( A1 => n140, A2 => n139, ZN => n219);
   U169 : NOR2_X1 port map( A1 => n246, A2 => n247, ZN => n239);
   U170 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => n246);
   U171 : NOR2_X1 port map( A1 => n190, A2 => n191, ZN => n183);
   U172 : NAND2_X1 port map( A1 => n93, A2 => n94, ZN => n87);
   U173 : AND2_X1 port map( A1 => n320, A2 => n319, ZN => n64);
   U174 : NAND2_X1 port map( A1 => n101, A2 => n102, ZN => n103);
   U175 : NAND2_X1 port map( A1 => n140, A2 => n305, ZN => n328);
   U176 : AND2_X1 port map( A1 => n196, A2 => n173, ZN => n188);
   U177 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => n196);
   U178 : INV_X1 port map( A => n267, ZN => n288);
   U179 : NAND2_X1 port map( A1 => n221, A2 => n222, ZN => n155);
   U180 : AOI21_X1 port map( B1 => n228, B2 => n229, A => n230, ZN => n221);
   U181 : NAND2_X1 port map( A1 => n58, A2 => n223, ZN => n222);
   U182 : INV_X1 port map( A => n231, ZN => n230);
   U183 : AND2_X1 port map( A1 => n227, A2 => n226, ZN => n228);
   U184 : INV_X1 port map( A => n124, ZN => n123);
   U185 : AND2_X1 port map( A1 => n269, A2 => n262, ZN => n65);
   U186 : XNOR2_X1 port map( A => n146, B => n108, ZN => DIFF(2));
   U187 : INV_X1 port map( A => B(28), ZN => n175);
   U188 : NAND2_X1 port map( A1 => A(24), A2 => n203, ZN => n172);
   U189 : INV_X1 port map( A => B(24), ZN => n203);
   U190 : INV_X1 port map( A => A(16), ZN => n298);
   U191 : INV_X1 port map( A => B(29), ZN => n158);
   U192 : INV_X1 port map( A => B(26), ZN => n193);
   U193 : NAND2_X1 port map( A1 => A(16), A2 => n297, ZN => n267);
   U194 : NAND2_X1 port map( A1 => A(17), A2 => n293, ZN => n268);
   U195 : INV_X1 port map( A => B(25), ZN => n200);
   U196 : NAND2_X1 port map( A1 => B(26), A2 => n194, ZN => n166);
   U197 : INV_X1 port map( A => B(14), ZN => n345);
   U198 : INV_X1 port map( A => A(10), ZN => n407);
   U199 : NAND2_X1 port map( A1 => B(24), A2 => n204, ZN => n174);
   U200 : INV_X1 port map( A => A(24), ZN => n204);
   U201 : NAND2_X1 port map( A1 => n386, A2 => n385, ZN => n212);
   U202 : INV_X1 port map( A => B(27), ZN => n181);
   U203 : INV_X1 port map( A => B(21), ZN => n256);
   U204 : INV_X1 port map( A => B(12), ZN => n359);
   U205 : NAND2_X1 port map( A1 => A(23), A2 => n237, ZN => n231);
   U206 : INV_X1 port map( A => B(23), ZN => n237);
   U207 : INV_X1 port map( A => B(15), ZN => n334);
   U208 : NAND2_X1 port map( A1 => B(23), A2 => n238, ZN => n227);
   U209 : INV_X1 port map( A => A(23), ZN => n238);
   U210 : NAND2_X1 port map( A1 => B(14), A2 => n346, ZN => n306);
   U211 : NAND2_X1 port map( A1 => B(19), A2 => n280, ZN => n269);
   U212 : INV_X1 port map( A => A(30), ZN => n144);
   U213 : NAND2_X1 port map( A1 => B(29), A2 => n159, ZN => n131);
   U214 : NAND2_X1 port map( A1 => B(15), A2 => n333, ZN => n305);
   U215 : OAI211_X1 port map( C1 => n391, C2 => n392, A => n26, B => n393, ZN 
                           => n390);
   U216 : NAND2_X1 port map( A1 => B(28), A2 => n176, ZN => n154);
   U217 : NAND2_X1 port map( A1 => A(10), A2 => n406, ZN => n319);
   U218 : INV_X1 port map( A => B(9), ZN => n378);
   U219 : NAND2_X1 port map( A1 => B(27), A2 => n182, ZN => n167);
   U220 : NAND2_X1 port map( A1 => A(4), A2 => n403, ZN => n101);
   U221 : NAND2_X1 port map( A1 => A(30), A2 => n145, ZN => n124);
   U222 : NAND2_X1 port map( A1 => n261, A2 => n262, ZN => n223);
   U223 : AND2_X1 port map( A1 => n269, A2 => n270, ZN => n263);
   U224 : NAND2_X1 port map( A1 => B(12), A2 => n360, ZN => n322);
   U225 : XNOR2_X1 port map( A => n275, B => n150, ZN => DIFF(1));
   U226 : OR2_X1 port map( A1 => n66, A2 => n408, ZN => DIFF(0));
   U227 : NAND2_X1 port map( A1 => A(3), A2 => n388, ZN => n110);
   U228 : AND2_X1 port map( A1 => A(8), A2 => n405, ZN => n68);
   U229 : INV_X1 port map( A => B(19), ZN => n279);
   U230 : NAND2_X1 port map( A1 => n326, A2 => n327, ZN => n216);
   U231 : INV_X1 port map( A => A(4), ZN => n316);
   U232 : INV_X1 port map( A => A(3), ZN => n389);
   U233 : XOR2_X1 port map( A => B(31), B => A(31), Z => n69);
   U234 : INV_X1 port map( A => B(20), ZN => n273);
   U235 : NAND2_X1 port map( A1 => B(20), A2 => n274, ZN => n224);
   U236 : INV_X1 port map( A => B(18), ZN => n289);
   U237 : NAND2_X1 port map( A1 => B(18), A2 => n290, ZN => n270);
   U238 : NOR2_X1 port map( A1 => B(4), A2 => n316, ZN => n313);
   U239 : NAND2_X1 port map( A1 => B(4), A2 => n316, ZN => n102);
   U240 : INV_X1 port map( A => B(4), ZN => n403);
   U241 : NAND2_X1 port map( A1 => A(28), A2 => n175, ZN => n125);
   U242 : INV_X1 port map( A => A(28), ZN => n176);
   U243 : NAND2_X1 port map( A1 => n41, A2 => n96, ZN => n99);
   U244 : OAI211_X1 port map( C1 => n313, C2 => n314, A => n97, B => n9, ZN => 
                           n311);
   U245 : NAND2_X1 port map( A1 => n97, A2 => n91, ZN => n396);
   U246 : NAND2_X1 port map( A1 => A(29), A2 => n158, ZN => n128);
   U247 : INV_X1 port map( A => A(29), ZN => n159);
   U248 : NAND2_X1 port map( A1 => n27, A2 => n64, ZN => n355);
   U249 : AOI21_X1 port map( B1 => n64, B2 => n27, A => n321, ZN => n361);
   U250 : INV_X1 port map( A => B(17), ZN => n293);
   U251 : NAND2_X1 port map( A1 => B(16), A2 => n298, ZN => n271);
   U252 : INV_X1 port map( A => B(16), ZN => n297);
   U253 : NAND2_X1 port map( A1 => B(13), A2 => n350, ZN => n323);
   U254 : INV_X1 port map( A => B(13), ZN => n349);
   U255 : INV_X1 port map( A => A(21), ZN => n257);
   U256 : NAND2_X1 port map( A1 => A(21), A2 => n256, ZN => n234);
   U257 : INV_X1 port map( A => B(30), ZN => n145);
   U258 : NAND2_X1 port map( A1 => B(30), A2 => n144, ZN => n130);
   U259 : INV_X1 port map( A => A(20), ZN => n274);
   U260 : NAND2_X1 port map( A1 => A(20), A2 => n273, ZN => n232);
   U261 : XNOR2_X1 port map( A => n286, B => n285, ZN => DIFF(18));
   U262 : NAND2_X1 port map( A1 => B(17), A2 => n294, ZN => n272);
   U263 : INV_X1 port map( A => A(17), ZN => n294);
   U264 : INV_X1 port map( A => B(22), ZN => n249);
   U265 : NAND2_X1 port map( A1 => B(22), A2 => n250, ZN => n226);
   U266 : NAND2_X1 port map( A1 => A(27), A2 => n181, ZN => n165);
   U267 : INV_X1 port map( A => A(27), ZN => n182);
   U268 : XNOR2_X1 port map( A => n69, B => n111, ZN => DIFF(31));
   U269 : NAND2_X1 port map( A1 => A(26), A2 => n193, ZN => n170);
   U270 : INV_X1 port map( A => A(26), ZN => n194);
   U271 : NOR2_X1 port map( A1 => B(5), A2 => n315, ZN => n314);
   U272 : INV_X1 port map( A => B(5), ZN => n402);
   U273 : NAND2_X1 port map( A1 => B(5), A2 => n315, ZN => n97);
   U274 : NAND2_X1 port map( A1 => A(9), A2 => n378, ZN => n79);
   U275 : INV_X1 port map( A => B(7), ZN => n398);
   U276 : NAND2_X1 port map( A1 => B(7), A2 => n404, ZN => n93);
   U277 : NAND2_X1 port map( A1 => A(2), A2 => n74, ZN => n107);
   U278 : INV_X1 port map( A => A(2), ZN => n387);
   U279 : INV_X1 port map( A => B(11), ZN => n375);
   U280 : NAND2_X1 port map( A1 => B(11), A2 => n376, ZN => n356);
   U281 : NAND2_X1 port map( A1 => A(19), A2 => n279, ZN => n262);
   U282 : INV_X1 port map( A => A(19), ZN => n280);
   U283 : INV_X1 port map( A => A(8), ZN => n369);
   U284 : NAND2_X1 port map( A1 => A(25), A2 => n200, ZN => n171);
   U285 : INV_X1 port map( A => A(25), ZN => n201);
   U286 : INV_X1 port map( A => B(10), ZN => n406);
   U287 : NAND2_X1 port map( A1 => B(10), A2 => n407, ZN => n364);
   U288 : NAND2_X1 port map( A1 => A(18), A2 => n289, ZN => n266);
   U289 : INV_X1 port map( A => A(18), ZN => n290);
   U290 : NAND2_X1 port map( A1 => A(13), A2 => n349, ZN => n304);
   U291 : INV_X1 port map( A => A(13), ZN => n350);
   U292 : NAND2_X1 port map( A1 => A(15), A2 => n334, ZN => n140);
   U293 : INV_X1 port map( A => A(15), ZN => n333);
   U294 : INV_X1 port map( A => B(6), ZN => n397);
   U295 : NAND2_X1 port map( A1 => B(6), A2 => n399, ZN => n91);
   U296 : INV_X1 port map( A => A(22), ZN => n250);
   U297 : NAND2_X1 port map( A1 => A(22), A2 => n249, ZN => n235);
   U298 : INV_X1 port map( A => A(7), ZN => n404);
   U299 : NAND2_X1 port map( A1 => A(7), A2 => n398, ZN => n94);
   U300 : NAND2_X1 port map( A1 => n28, A2 => n32, ZN => n338);
   U301 : NOR2_X1 port map( A1 => n210, A2 => n211, ZN => n209);
   U302 : NOR2_X1 port map( A1 => n321, A2 => n210, ZN => n317);
   U303 : NAND4_X1 port map( A1 => n322, A2 => n323, A3 => n306, A4 => n305, ZN
                           => n210);
   U304 : NAND2_X1 port map( A1 => n359, A2 => A(12), ZN => n302);
   U305 : INV_X1 port map( A => A(12), ZN => n360);
   U306 : OAI21_X1 port map( B1 => n147, B2 => n217, A => n149, ZN => n108);
   U307 : NAND2_X1 port map( A1 => A(5), A2 => n402, ZN => n96);
   U308 : INV_X1 port map( A => A(5), ZN => n315);
   U309 : XNOR2_X1 port map( A => n6, B => n103, ZN => DIFF(4));
   U310 : NAND2_X1 port map( A1 => n86, A2 => n102, ZN => n100);
   U311 : OAI21_X1 port map( B1 => n372, B2 => n373, A => n319, ZN => n371);
   U312 : XNOR2_X1 port map( A => n152, B => n151, ZN => DIFF(29));
   U313 : NAND2_X1 port map( A1 => n109, A2 => n110, ZN => n104);
   U314 : OAI21_X1 port map( B1 => n73, B2 => n387, A => n110, ZN => n386);
   U315 : NAND2_X1 port map( A1 => B(3), A2 => n389, ZN => n385);
   U316 : NAND2_X1 port map( A1 => B(3), A2 => n389, ZN => n109);
   U317 : INV_X1 port map( A => B(3), ZN => n388);
   U318 : NAND2_X1 port map( A1 => A(14), A2 => n345, ZN => n303);
   U319 : INV_X1 port map( A => A(14), ZN => n346);
   U320 : INV_X1 port map( A => A(9), ZN => n368);
   U321 : NAND2_X1 port map( A1 => B(9), A2 => n368, ZN => n365);
   U322 : NAND4_X1 port map( A1 => n356, A2 => n364, A3 => n365, A4 => n81, ZN 
                           => n211);
   U323 : NAND2_X1 port map( A1 => n25, A2 => n71, ZN => n276);
   U324 : NOR2_X1 port map( A1 => B(0), A2 => n394, ZN => n391);
   U325 : NAND2_X1 port map( A1 => A(0), A2 => n71, ZN => n327);
   U326 : INV_X1 port map( A => A(0), ZN => n394);
   U327 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => n88);
   U328 : NAND2_X1 port map( A1 => n277, A2 => n149, ZN => n275);
   U329 : INV_X1 port map( A => B(8), ZN => n405);
   U330 : NOR2_X1 port map( A1 => B(8), A2 => n369, ZN => n366);
   U331 : NAND2_X1 port map( A1 => B(8), A2 => n369, ZN => n81);
   U332 : AND2_X1 port map( A1 => n220, A2 => n70, ZN => n299);
   U333 : AND2_X1 port map( A1 => n139, A2 => n140, ZN => n70);
   U334 : INV_X1 port map( A => A(11), ZN => n376);
   U335 : NAND2_X1 port map( A1 => n20, A2 => n375, ZN => n320);
   U336 : AOI21_X1 port map( B1 => n195, B2 => n61, A => n188, ZN => n192);
   U337 : XNOR2_X1 port map( A => n99, B => n98, ZN => DIFF(5));
   U338 : AND2_X1 port map( A1 => n382, A2 => n385, ZN => n393);
   U339 : NAND2_X1 port map( A1 => n26, A2 => n382, ZN => n325);
   U340 : NAND2_X1 port map( A1 => n18, A2 => n92, ZN => n90);
   U341 : NAND2_X1 port map( A1 => n382, A2 => n107, ZN => n146);
   U342 : AOI21_X1 port map( B1 => n251, B2 => n225, A => n244, ZN => n248);
   U343 : AOI21_X1 port map( B1 => n47, B2 => n6, A => n33, ZN => n83);
   U344 : NAND2_X1 port map( A1 => n47, A2 => n86, ZN => n357);
   U345 : NAND2_X1 port map( A1 => n47, A2 => n6, ZN => n363);
   U346 : NAND4_X1 port map( A1 => n337, A2 => n47, A3 => n323, A4 => n6, ZN =>
                           n336);
   U347 : NAND4_X1 port map( A1 => n38, A2 => n40, A3 => n28, A4 => n47, ZN => 
                           n220);
   U348 : NAND2_X1 port map( A1 => A(6), A2 => n397, ZN => n89);
   U349 : INV_X1 port map( A => A(6), ZN => n399);
   U350 : XNOR2_X1 port map( A => n278, B => n65, ZN => DIFF(19));
   U351 : XNOR2_X1 port map( A => n10, B => n296, ZN => DIFF(16));
   U352 : NOR2_X1 port map( A1 => n281, A2 => n282, ZN => n278);
   U353 : AOI21_X1 port map( B1 => n10, B2 => n239, A => n240, ZN => n236);
   U354 : AOI21_X1 port map( B1 => n10, B2 => n183, A => n184, ZN => n177);
   U355 : NAND2_X1 port map( A1 => n52, A2 => n271, ZN => n295);
   U356 : OAI211_X1 port map( C1 => n10, C2 => n288, A => n271, B => n272, ZN 
                           => n287);
   U357 : NAND2_X1 port map( A1 => n82, A2 => n363, ZN => n80);
   U358 : NAND2_X1 port map( A1 => n381, A2 => n357, ZN => n380);
   U359 : NOR2_X1 port map( A1 => B(1), A2 => n21, ZN => n392);
   U360 : NAND2_X1 port map( A1 => B(1), A2 => n384, ZN => n218);
   U361 : NAND2_X1 port map( A1 => B(1), A2 => n384, ZN => n277);
   U362 : INV_X1 port map( A => B(1), ZN => n72);
   U363 : OAI21_X1 port map( B1 => n44, B2 => n49, A => n96, ZN => n92);
   U364 : XNOR2_X1 port map( A => n87, B => n88, ZN => DIFF(7));
   U365 : OAI21_X1 port map( B1 => n247, B2 => n34, A => n241, ZN => n253);
   U366 : OAI21_X1 port map( B1 => n48, B2 => n255, A => n260, ZN => n259);
   U367 : OAI211_X1 port map( C1 => n117, C2 => n34, A => n121, B => n63, ZN =>
                           n152);
   U368 : OAI21_X1 port map( B1 => n34, B2 => n247, A => n241, ZN => n251);
   U369 : OAI21_X1 port map( B1 => n48, B2 => n191, A => n185, ZN => n195);
   U370 : AOI21_X1 port map( B1 => n48, B2 => n267, A => n284, ZN => n281);
   U371 : NAND2_X1 port map( A1 => n31, A2 => n72, ZN => n149);
   U372 : NAND2_X1 port map( A1 => n31, A2 => n72, ZN => n326);
   U373 : INV_X1 port map( A => A(1), ZN => n384);
   U374 : INV_X1 port map( A => B(0), ZN => n71);
   U375 : INV_X1 port map( A => n74, ZN => n73);
   U376 : INV_X1 port map( A => B(2), ZN => n74);
   U377 : NOR2_X1 port map( A1 => n77, A2 => n78, ZN => n76);
   U378 : INV_X1 port map( A => n79, ZN => n77);
   U379 : NOR2_X1 port map( A1 => n68, A2 => n85, ZN => n84);
   U380 : XNOR2_X1 port map( A => n95, B => n92, ZN => DIFF(6));
   U381 : XNOR2_X1 port map( A => n104, B => n105, ZN => DIFF(3));
   U382 : OAI21_X1 port map( B1 => n106, B2 => n46, A => n107, ZN => n105);
   U383 : INV_X1 port map( A => n108, ZN => n106);
   U384 : NAND3_X1 port map( A1 => n52, A2 => n116, A3 => n120, ZN => n115);
   U385 : INV_X1 port map( A => n131, ZN => n134);
   U386 : INV_X1 port map( A => n150, ZN => n147);
   U387 : XNOR2_X1 port map( A => n161, B => n160, ZN => DIFF(28));
   U388 : INV_X1 port map( A => n153, ZN => n162);
   U389 : NOR2_X1 port map( A1 => n179, A2 => n180, ZN => n178);
   U390 : INV_X1 port map( A => n165, ZN => n180);
   U391 : INV_X1 port map( A => n167, ZN => n179);
   U392 : INV_X1 port map( A => n170, ZN => n189);
   U393 : NAND2_X1 port map( A1 => n61, A2 => n166, ZN => n186);
   U394 : NAND2_X1 port map( A1 => n61, A2 => n166, ZN => n190);
   U395 : XNOR2_X1 port map( A => n197, B => n198, ZN => DIFF(25));
   U396 : INV_X1 port map( A => n174, ZN => n199);
   U397 : OAI21_X1 port map( B1 => n206, B2 => n207, A => n156, ZN => n205);
   U398 : INV_X1 port map( A => n191, ZN => n156);
   U399 : NAND3_X1 port map( A1 => n143, A2 => n39, A3 => n141, ZN => n207);
   U400 : NAND3_X1 port map( A1 => n208, A2 => n47, A3 => n8, ZN => n143);
   U401 : INV_X1 port map( A => n109, ZN => n214);
   U402 : NOR2_X1 port map( A1 => n46, A2 => n217, ZN => n215);
   U403 : INV_X1 port map( A => n277, ZN => n217);
   U404 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => n206);
   U405 : INV_X1 port map( A => n155, ZN => n185);
   U406 : INV_X1 port map( A => n235, ZN => n245);
   U407 : INV_X1 port map( A => n234, ZN => n244);
   U408 : XNOR2_X1 port map( A => n252, B => n253, ZN => DIFF(21));
   U409 : INV_X1 port map( A => n232, ZN => n254);
   U410 : XNOR2_X1 port map( A => n258, B => n259, ZN => DIFF(20));
   U411 : INV_X1 port map( A => n223, ZN => n260);
   U412 : NAND3_X1 port map( A1 => n263, A2 => n264, A3 => n265, ZN => n261);
   U413 : NAND3_X1 port map( A1 => n267, A2 => n268, A3 => n266, ZN => n264);
   U414 : INV_X1 port map( A => n29, ZN => n283);
   U415 : NAND3_X1 port map( A1 => n271, A2 => n29, A3 => n272, ZN => n284);
   U416 : NAND3_X1 port map( A1 => n319, A2 => n320, A3 => n35, ZN => n318);
   U417 : XNOR2_X1 port map( A => n328, B => n329, ZN => DIFF(15));
   U418 : INV_X1 port map( A => n306, ZN => n331);
   U419 : INV_X1 port map( A => n332, ZN => n330);
   U420 : NAND3_X1 port map( A1 => n335, A2 => n304, A3 => n336, ZN => n332);
   U421 : INV_X1 port map( A => n338, ZN => n337);
   U422 : NAND2_X1 port map( A1 => n343, A2 => n344, ZN => n342);
   U423 : NOR2_X1 port map( A1 => n30, A2 => n312, ZN => n343);
   U424 : INV_X1 port map( A => n93, ZN => n312);
   U425 : NOR2_X1 port map( A1 => n30, A2 => n37, ZN => n339);
   U426 : INV_X1 port map( A => n340, ZN => n353);
   U427 : INV_X1 port map( A => n356, ZN => n321);
   U428 : XNOR2_X1 port map( A => n370, B => n371, ZN => DIFF(11));
   U429 : INV_X1 port map( A => n19, ZN => n373);
   U430 : INV_X1 port map( A => n374, ZN => n372);
   U431 : NAND3_X1 port map( A1 => n14, A2 => n385, A3 => n382, ZN => n307);
   U432 : NOR2_X1 port map( A1 => n148, A2 => n66, ZN => n383);
   U433 : INV_X1 port map( A => n218, ZN => n148);
   U434 : NOR2_X1 port map( A1 => n68, A2 => n33, ZN => n381);
   U435 : NOR2_X1 port map( A1 => n400, A2 => n401, ZN => n395);
   U436 : INV_X1 port map( A => n96, ZN => n401);
   U437 : INV_X1 port map( A => n101, ZN => n400);
   U438 : NOR2_X1 port map( A1 => n85, A2 => n78, ZN => n379);
   U439 : INV_X1 port map( A => n17, ZN => n78);
   U440 : INV_X1 port map( A => n22, ZN => n85);
   U441 : INV_X1 port map( A => n276, ZN => n408);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BARREL_SHIFTER_N32 is

   port( CONF : in std_logic;  DATA1, DATA2 : in std_logic_vector (31 downto 0)
         ;  OUTPUT : out std_logic_vector (31 downto 0));

end BARREL_SHIFTER_N32;

architecture SYN_BEHAVIOR of BARREL_SHIFTER_N32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal net46810, net46815, net46817, net46819, net46838, net46850, net46851,
      net46854, net46856, net46857, net46859, net46877, net46878, net46879, 
      net46880, net46881, net46901, net46911, net46934, net46936, net46949, 
      net46956, net46957, net46966, net46967, net46971, net46972, net46973, 
      net46974, net46975, net46978, net46980, net46988, net46991, net46993, 
      net46994, net46995, net47004, net47009, net47010, net47012, net47013, 
      net47018, net47019, net47025, net47026, net47028, net47037, net47039, 
      net47042, net47043, net47049, net47050, net47060, net47065, net47109, 
      net47150, net47157, net47177, net47178, net47183, net47184, net47187, 
      net47197, net50841, net50839, net50837, net50835, net50833, net50831, 
      net50827, net50871, net50869, net50867, net50865, net50863, net50861, 
      net50857, net50905, net50901, net50899, net50897, net50895, net50893, 
      net50891, net50889, net51555, net51553, net51551, net51549, net51547, 
      net51543, net51599, net51703, net51702, net52169, net52168, net52292, 
      net54951, net54952, net55100, net55209, net55611, net55654, net55672, 
      net55714, net55741, net55740, net55739, net55767, net55782, net55789, 
      net55829, net55828, net55852, net55902, net55928, net55953, net55980, 
      net55991, net56027, net56098, net56118, net56120, net56146, net56178, 
      net56183, net56186, net56192, net56195, net56207, net56216, net56225, 
      net56256, net56277, net56276, net56281, net56284, net51559, net46816, 
      net55634, net50903, net46998, net56159, net51557, net54992, net51541, 
      net46981, net46818, net47003, net46958, net47038, net47014, net47002, 
      net47000, net46999, net46979, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
      n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
      n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
      n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
      n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
      n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
      n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
      n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
      n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
      n338, n339, n340 : std_logic;

begin
   
   U2 : MUX2_X1 port map( A => net46859, B => net46911, S => net50839, Z => 
                           n262);
   U3 : INV_X1 port map( A => net50837, ZN => net50835);
   U4 : BUF_X1 port map( A => net55767, Z => n1);
   U5 : CLKBUF_X1 port map( A => DATA2(4), Z => net55767);
   U6 : CLKBUF_X1 port map( A => net55828, Z => n2);
   U7 : MUX2_X1 port map( A => n15, B => net47026, S => net50871, Z => net47013
                           );
   U8 : CLKBUF_X1 port map( A => net46859, Z => net55902);
   U9 : MUX2_X1 port map( A => n54, B => n55, S => net50839, Z => n61);
   U10 : INV_X1 port map( A => net50837, ZN => net50827);
   U11 : AND2_X1 port map( A1 => net55902, A2 => net50841, ZN => n3);
   U12 : INV_X2 port map( A => DATA2(2), ZN => net50841);
   U13 : MUX2_X1 port map( A => n123, B => net47157, S => net50837, Z => n85);
   U14 : MUX2_X1 port map( A => n274, B => n252, S => net50871, Z => n264);
   U15 : MUX2_X1 port map( A => net47013, B => net47025, S => net50905, Z => 
                           n198);
   U16 : MUX2_X1 port map( A => net46981, B => net47028, S => net50839, Z => 
                           n17);
   U17 : MUX2_X1 port map( A => n33, B => n291, S => DATA2(2), Z => n251);
   U18 : INV_X1 port map( A => net51557, ZN => n4);
   U19 : MUX2_X2 port map( A => n274, B => n292, S => net50865, Z => n285);
   U20 : OR2_X1 port map( A1 => net55829, A2 => net46973, ZN => n5);
   U21 : OR2_X1 port map( A1 => net51703, A2 => net46879, ZN => n6);
   U22 : NAND3_X1 port map( A1 => n5, A2 => n6, A3 => net47065, ZN => net47003)
                           ;
   U23 : AND2_X1 port map( A1 => net51555, A2 => net54952, ZN => n7);
   U24 : INV_X2 port map( A => n7, ZN => n66);
   U25 : MUX2_X1 port map( A => net47003, B => net47050, S => net50839, Z => 
                           net47049);
   U26 : MUX2_X1 port map( A => n233, B => n273, S => net50835, Z => n234);
   U27 : INV_X2 port map( A => DATA2(2), ZN => net50837);
   U28 : MUX2_X1 port map( A => n264, B => n275, S => net50899, Z => n265);
   U29 : BUF_X2 port map( A => net46816, Z => net51599);
   U30 : INV_X1 port map( A => n8, ZN => net46878);
   U31 : MUX2_X1 port map( A => n61, B => n78, S => net50863, Z => n70);
   U32 : INV_X1 port map( A => net50867, ZN => net50863);
   U33 : INV_X1 port map( A => net50869, ZN => net50857);
   U34 : MUX2_X1 port map( A => n40, B => n323, S => net50839, Z => n325);
   U35 : MUX2_X1 port map( A => n327, B => n304, S => net50867, Z => net46838);
   U36 : INV_X2 port map( A => net50867, ZN => net50865);
   U37 : MUX2_X1 port map( A => n113, B => n154, S => DATA2(2), Z => n114);
   U38 : AND2_X2 port map( A1 => net54952, A2 => net55714, ZN => n8);
   U39 : INV_X1 port map( A => net50841, ZN => n9);
   U40 : CLKBUF_X1 port map( A => n4, Z => net52169);
   U41 : MUX2_X1 port map( A => net46967, B => n235, S => net50863, Z => n227);
   U42 : BUF_X2 port map( A => net46818, Z => n10);
   U43 : AND2_X1 port map( A1 => net51555, A2 => net54951, ZN => net55672);
   U44 : CLKBUF_X1 port map( A => net51553, Z => net51551);
   U45 : AND2_X2 port map( A1 => net51553, A2 => net55953, ZN => net55611);
   U46 : INV_X1 port map( A => net56183, ZN => n11);
   U47 : MUX2_X1 port map( A => n264, B => n253, S => net50905, Z => n254);
   U48 : MUX2_X1 port map( A => n30, B => net46936, S => net50841, Z => n244);
   U49 : MUX2_X1 port map( A => n245, B => n236, S => net50905, Z => n237);
   U50 : BUF_X2 port map( A => net46816, Z => net56118);
   U51 : INV_X1 port map( A => net56183, ZN => n12);
   U52 : MUX2_X2 port map( A => n311, B => n312, S => net50839, Z => n333);
   U53 : MUX2_X1 port map( A => n326, B => n335, S => net50905, Z => n330);
   U54 : NOR2_X1 port map( A1 => DATA2(4), A2 => net55782, ZN => net54992);
   U55 : AND2_X2 port map( A1 => net51555, A2 => n31, ZN => n32);
   U56 : NAND2_X2 port map( A1 => net55714, A2 => n31, ZN => net55829);
   U57 : OR2_X2 port map( A1 => net47009, A2 => net51557, ZN => net56183);
   U58 : MUX2_X1 port map( A => n96, B => n87, S => net50905, Z => n88);
   U59 : INV_X1 port map( A => net50903, ZN => net50889);
   U60 : MUX2_X1 port map( A => n313, B => n289, S => net50861, Z => n303);
   U61 : INV_X1 port map( A => net50867, ZN => net50861);
   U62 : MUX2_X1 port map( A => n13, B => net47000, S => net50905, Z => 
                           net46999);
   U63 : OAI22_X1 port map( A1 => net51549, A2 => net46998, B1 => net46999, B2 
                           => net51543, ZN => OUTPUT(16));
   U64 : INV_X2 port map( A => DATA2(0), ZN => net50905);
   U65 : MUX2_X1 port map( A => net46979, B => n15, S => net50871, Z => n13);
   U66 : MUX2_X1 port map( A => n13, B => net46978, S => net50893, Z => 
                           net46988);
   U67 : INV_X2 port map( A => DATA2(1), ZN => net50871);
   U68 : INV_X1 port map( A => n17, ZN => n15);
   U69 : INV_X2 port map( A => DATA2(2), ZN => net50839);
   U70 : INV_X1 port map( A => net47002, ZN => net46979);
   U71 : MUX2_X1 port map( A => net46979, B => net46956, S => net50863, Z => 
                           net46966);
   U72 : MUX2_X1 port map( A => net47003, B => net46958, S => net50831, Z => 
                           net47002);
   U73 : INV_X1 port map( A => net50837, ZN => net50831);
   U74 : MUX2_X1 port map( A => n14, B => net47014, S => net50867, Z => 
                           net47000);
   U75 : MUX2_X1 port map( A => net47013, B => net47000, S => net50893, Z => 
                           net47012);
   U76 : INV_X1 port map( A => DATA2(1), ZN => net50867);
   U77 : INV_X1 port map( A => net47038, ZN => net47014);
   U78 : MUX2_X1 port map( A => net47037, B => net47014, S => DATA2(1), Z => 
                           net47025);
   U79 : MUX2_X1 port map( A => net55789, B => net47039, S => net50841, Z => 
                           net47038);
   U80 : INV_X1 port map( A => n16, ZN => n14);
   U81 : MUX2_X1 port map( A => net46967, B => n14, S => net50871, Z => 
                           net46978);
   U82 : MUX2_X1 port map( A => net56195, B => net56192, S => net50839, Z => 
                           n16);
   U83 : INV_X1 port map( A => DATA2(0), ZN => net50901);
   U84 : INV_X1 port map( A => DATA2(0), ZN => net50903);
   U85 : INV_X1 port map( A => DATA2(1), ZN => net50869);
   U86 : MUX2_X1 port map( A => net46936, B => net46981, S => net50839, Z => 
                           net46980);
   U87 : MUX2_X1 port map( A => net46981, B => net47028, S => net50831, Z => 
                           net47042);
   U88 : INV_X1 port map( A => DATA1(3), ZN => net46879);
   U89 : BUF_X2 port map( A => net56159, Z => net51702);
   U90 : INV_X1 port map( A => DATA1(11), ZN => net46973);
   U91 : OAI221_X1 port map( B1 => net51702, B2 => n20, C1 => net56118, C2 => 
                           n18, A => n21, ZN => net46958);
   U92 : MUX2_X1 port map( A => net46911, B => net46958, S => net50841, Z => 
                           net46957);
   U93 : MUX2_X1 port map( A => net46958, B => net56186, S => net50831, Z => 
                           net47019);
   U94 : MUX2_X1 port map( A => net46911, B => net46958, S => net50833, Z => 
                           net46972);
   U95 : AOI22_X1 port map( A1 => net55611, A2 => DATA1(31), B1 => net56216, B2
                           => DATA1(23), ZN => n21);
   U96 : INV_X1 port map( A => DATA1(15), ZN => n18);
   U97 : OAI221_X1 port map( B1 => net51702, B2 => n18, C1 => net51599, C2 => 
                           net46819, A => n19, ZN => net46859);
   U98 : INV_X1 port map( A => DATA1(7), ZN => n20);
   U99 : OAI221_X1 port map( B1 => net55828, B2 => n20, C1 => net46819, C2 => 
                           net52292, A => n22, ZN => net47050);
   U100 : OAI221_X1 port map( B1 => net55829, B2 => net46973, C1 => net56207, 
                           C2 => net46879, A => net47065, ZN => net56186);
   U101 : AOI22_X1 port map( A1 => net55741, A2 => DATA1(3), B1 => net56216, B2
                           => DATA1(27), ZN => net46975);
   U102 : INV_X1 port map( A => net56159, ZN => net46881);
   U103 : AOI22_X1 port map( A1 => DATA1(19), A2 => net46881, B1 => net55739, 
                           B2 => DATA1(11), ZN => net46880);
   U104 : AOI22_X1 port map( A1 => net55740, A2 => DATA1(7), B1 => net56178, B2
                           => DATA1(31), ZN => n19);
   U105 : AOI22_X1 port map( A1 => DATA1(15), A2 => net56178, B1 => net55672, 
                           B2 => DATA1(31), ZN => n22);
   U106 : INV_X1 port map( A => DATA1(31), ZN => net46817);
   U107 : INV_X1 port map( A => DATA1(23), ZN => net46819);
   U108 : AOI22_X1 port map( A1 => net56281, A2 => DATA1(23), B1 => net55611, 
                           B2 => DATA1(15), ZN => net47178);
   U109 : AOI221_X1 port map( B1 => DATA1(7), B2 => n8, C1 => DATA1(15), C2 => 
                           net56098, A => net46815, ZN => net46810);
   U110 : OAI221_X1 port map( B1 => net47043, B2 => n10, C1 => net55654, C2 => 
                           n23, A => n24, ZN => net46981);
   U111 : MUX2_X1 port map( A => net46936, B => net46981, S => net50831, Z => 
                           net46995);
   U112 : AOI22_X1 port map( A1 => n37, A2 => DATA1(29), B1 => net56216, B2 => 
                           DATA1(21), ZN => n24);
   U113 : INV_X1 port map( A => DATA1(13), ZN => n23);
   U114 : OR2_X1 port map( A1 => net51703, A2 => n23, ZN => net55928);
   U115 : OAI222_X1 port map( A1 => net47043, A2 => net56276, B1 => net47184, 
                           B2 => net52169, C1 => n23, C2 => net47109, ZN => 
                           net47157);
   U116 : BUF_X2 port map( A => net46818, Z => net51703);
   U117 : NAND2_X1 port map( A1 => net51541, A2 => net54992, ZN => net46818);
   U118 : INV_X1 port map( A => net51557, ZN => net51541);
   U119 : NAND2_X1 port map( A1 => net51541, A2 => net54992, ZN => net56159);
   U120 : BUF_X1 port map( A => CONF, Z => net51557);
   U121 : CLKBUF_X1 port map( A => DATA2(3), Z => n25);
   U122 : AND2_X1 port map( A1 => net55767, A2 => n25, ZN => net54952);
   U123 : INV_X1 port map( A => DATA2(4), ZN => net47187);
   U124 : INV_X1 port map( A => DATA2(3), ZN => net47010);
   U125 : INV_X1 port map( A => DATA2(3), ZN => net55782);
   U126 : BUF_X1 port map( A => DATA2(3), Z => net56120);
   U127 : CLKBUF_X1 port map( A => DATA2(4), Z => net55980);
   U128 : INV_X2 port map( A => net51557, ZN => net55714);
   U129 : BUF_X1 port map( A => CONF, Z => net51559);
   U130 : INV_X2 port map( A => net51547, ZN => net51543);
   U131 : BUF_X2 port map( A => net55634, Z => net51547);
   U132 : INV_X1 port map( A => n4, ZN => net55634);
   U133 : NAND2_X1 port map( A1 => net56225, A2 => net55634, ZN => net47197);
   U134 : BUF_X1 port map( A => net55634, Z => net51549);
   U135 : MUX2_X1 port map( A => net46993, B => net47004, S => net50893, Z => 
                           net46998);
   U136 : INV_X1 port map( A => net50903, ZN => net50893);
   U137 : MUX2_X1 port map( A => net46838, B => net46857, S => net50903, Z => 
                           net46856);
   U138 : INV_X1 port map( A => net50903, ZN => net50891);
   U139 : CLKBUF_X3 port map( A => net51559, Z => net51553);
   U140 : BUF_X2 port map( A => net51559, Z => net51555);
   U141 : AND2_X2 port map( A1 => net51555, A2 => net55209, ZN => net56216);
   U142 : NAND2_X1 port map( A1 => net55100, A2 => net55714, ZN => net46816);
   U143 : NAND3_X1 port map( A1 => net55991, A2 => DATA1(7), A3 => net51553, ZN
                           => net47177);
   U144 : MUX2_X1 port map( A => n236, B => n227, S => net50905, Z => n228);
   U145 : MUX2_X1 port map( A => net46934, B => n263, S => net50861, Z => n253)
                           ;
   U146 : CLKBUF_X1 port map( A => net51702, Z => net56284);
   U147 : AND2_X1 port map( A1 => net51555, A2 => net54951, ZN => net56281);
   U148 : BUF_X1 port map( A => net47150, Z => net56276);
   U149 : BUF_X1 port map( A => net47150, Z => net56277);
   U150 : BUF_X1 port map( A => n123, Z => n26);
   U151 : INV_X1 port map( A => net51547, ZN => net56256);
   U152 : CLKBUF_X1 port map( A => n7, Z => n27);
   U153 : BUF_X1 port map( A => net54951, Z => net56225);
   U154 : AND2_X1 port map( A1 => net55767, A2 => net47010, ZN => net54951);
   U155 : AND2_X2 port map( A1 => net51553, A2 => net55953, ZN => n37);
   U156 : MUX2_X1 port map( A => n184, B => net47026, S => net50861, Z => n190)
                           ;
   U157 : AND2_X1 port map( A1 => net47187, A2 => net47010, ZN => net55209);
   U158 : CLKBUF_X1 port map( A => net51702, Z => net56207);
   U159 : AOI221_X1 port map( B1 => net55852, B2 => DATA1(16), C1 => n27, C2 =>
                           DATA1(24), A => n52, ZN => n55);
   U160 : BUF_X1 port map( A => n143, Z => n28);
   U161 : OAI221_X1 port map( B1 => n194, B2 => net51703, C1 => net56118, C2 =>
                           n240, A => n193, ZN => net56195);
   U162 : OAI221_X1 port map( B1 => net55829, B2 => n212, C1 => net51702, C2 =>
                           n161, A => n160, ZN => net56192);
   U163 : MUX2_X1 port map( A => n249, B => n271, S => net50871, Z => n261);
   U164 : AND2_X1 port map( A1 => net55209, A2 => net51555, ZN => net56178);
   U165 : OAI211_X1 port map( C1 => net46901, C2 => n269, A => n267, B => n268,
                           ZN => n29);
   U166 : NAND3_X1 port map( A1 => n34, A2 => net55928, A3 => n230, ZN => n30);
   U167 : INV_X1 port map( A => net46881, ZN => net56146);
   U168 : AND2_X1 port map( A1 => net47187, A2 => net47010, ZN => n31);
   U169 : CLKBUF_X1 port map( A => n11, Z => net56098);
   U170 : MUX2_X1 port map( A => n69, B => n86, S => net50857, Z => n79);
   U171 : OAI221_X1 port map( B1 => n212, B2 => net51703, C1 => net51599, C2 =>
                           n280, A => n211, ZN => n33);
   U172 : INV_X1 port map( A => n1, ZN => net56027);
   U173 : MUX2_X1 port map( A => n206, B => n214, S => net50871, Z => net46993)
                           ;
   U174 : MUX2_X1 port map( A => net56195, B => n33, S => n9, Z => n219);
   U175 : MUX2_X1 port map( A => net47037, B => n175, S => net50869, Z => n185)
                           ;
   U176 : CLKBUF_X1 port map( A => net55100, Z => net55991);
   U177 : AND2_X1 port map( A1 => net47187, A2 => net56120, ZN => net55953);
   U178 : CLKBUF_X1 port map( A => n4, Z => net52168);
   U179 : AND2_X1 port map( A1 => net47187, A2 => net47010, ZN => net55100);
   U180 : OR2_X1 port map( A1 => net55829, A2 => net46851, ZN => n34);
   U181 : MUX2_X1 port map( A => n190, B => n185, S => net50901, Z => n186);
   U182 : MUX2_X1 port map( A => n253, B => n245, S => net50905, Z => n246);
   U183 : MUX2_X1 port map( A => n190, B => net47025, S => net50899, Z => n191)
                           ;
   U184 : MUX2_X1 port map( A => net46966, B => net46978, S => net50905, Z => 
                           n216);
   U185 : INV_X1 port map( A => net50901, ZN => net50895);
   U186 : MUX2_X1 port map( A => n293, B => n285, S => net50905, Z => n286);
   U187 : INV_X1 port map( A => net50901, ZN => net50897);
   U188 : MUX2_X1 port map( A => n333, B => n313, S => net50865, Z => n35);
   U189 : MUX2_X1 port map( A => n284, B => n263, S => net50871, Z => n275);
   U190 : MUX2_X1 port map( A => n175, B => n156, S => net50871, Z => n168);
   U191 : BUF_X1 port map( A => n291, Z => n36);
   U192 : INV_X1 port map( A => net47197, ZN => net55852);
   U193 : INV_X1 port map( A => net56183, ZN => net55741);
   U194 : MUX2_X1 port map( A => n125, B => n105, S => net50869, Z => n116);
   U195 : MUX2_X1 port map( A => n103, B => n143, S => n9, Z => n104);
   U196 : NAND2_X1 port map( A1 => n4, A2 => n31, ZN => net55828);
   U197 : NAND2_X1 port map( A1 => net55100, A2 => n4, ZN => net55654);
   U198 : OR2_X1 port map( A1 => net55654, A2 => n139, ZN => n38);
   U199 : OR2_X1 port map( A1 => n204, A2 => net47109, ZN => n39);
   U200 : NAND3_X1 port map( A1 => n38, A2 => n39, A3 => n49, ZN => n113);
   U201 : NAND2_X1 port map( A1 => net51555, A2 => net55209, ZN => net47150);
   U202 : MUX2_X1 port map( A => n156, B => n134, S => net50869, Z => n146);
   U203 : MUX2_X1 port map( A => n176, B => n168, S => net50905, Z => n169);
   U204 : MUX2_X1 port map( A => net46934, B => net46956, S => net50867, Z => 
                           n236);
   U205 : OAI221_X1 port map( B1 => net56146, B2 => n180, C1 => net56118, C2 =>
                           n223, A => n179, ZN => net55789);
   U206 : MUX2_X1 port map( A => n134, B => n115, S => net50871, Z => n126);
   U207 : MUX2_X1 port map( A => n87, B => n79, S => net50905, Z => n80);
   U208 : MUX2_X1 port map( A => n252, B => n235, S => net50871, Z => n245);
   U209 : AND3_X1 port map( A1 => n41, A2 => n42, A3 => n278, ZN => n40);
   U210 : OR2_X1 port map( A1 => net51702, A2 => n280, ZN => n41);
   U211 : OR2_X1 port map( A1 => net55654, A2 => n279, ZN => n42);
   U212 : NAND3_X1 port map( A1 => n41, A2 => n42, A3 => n278, ZN => n322);
   U213 : INV_X1 port map( A => net56183, ZN => net55739);
   U214 : INV_X1 port map( A => net56183, ZN => net55740);
   U215 : MUX2_X1 port map( A => n157, B => n146, S => net50905, Z => n147);
   U216 : MUX2_X1 port map( A => n135, B => n126, S => net50905, Z => n127);
   U217 : MUX2_X1 port map( A => n167, B => n145, S => net50871, Z => n157);
   U218 : MUX2_X1 port map( A => n116, B => n106, S => net50905, Z => n107);
   U219 : NAND3_X1 port map( A1 => n44, A2 => n45, A3 => n82, ZN => n43);
   U220 : OR2_X1 port map( A1 => net55654, A2 => n161, ZN => n44);
   U221 : OR2_X1 port map( A1 => net47150, A2 => n212, ZN => n45);
   U222 : NAND3_X1 port map( A1 => n44, A2 => n45, A3 => n82, ZN => n132);
   U223 : MUX2_X1 port map( A => n105, B => n86, S => net50869, Z => n96);
   U224 : MUX2_X1 port map( A => n95, B => n78, S => net50871, Z => n87);
   U225 : NAND3_X1 port map( A1 => n48, A2 => n47, A3 => n138, ZN => n46);
   U226 : AOI221_X1 port map( B1 => net55852, B2 => DATA1(17), C1 => n27, C2 =>
                           DATA1(25), A => n62, ZN => n64);
   U227 : OAI221_X1 port map( B1 => n298, B2 => net51702, C1 => n2, C2 => n297,
                           A => n296, ZN => n300);
   U228 : OR2_X1 port map( A1 => n10, A2 => n139, ZN => n47);
   U229 : OR2_X1 port map( A1 => net55654, A2 => n258, ZN => n48);
   U230 : NAND3_X1 port map( A1 => n48, A2 => n47, A3 => n138, ZN => net47039);
   U231 : INV_X1 port map( A => n12, ZN => net46901);
   U232 : INV_X1 port map( A => net50837, ZN => net50833);
   U233 : NOR2_X1 port map( A1 => net46851, A2 => net51702, ZN => n309);
   U234 : AOI211_X1 port map( C1 => n310, C2 => net52169, A => n309, B => n308,
                           ZN => n312);
   U235 : INV_X1 port map( A => n29, ZN => n311);
   U236 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => n310);
   U237 : NAND2_X1 port map( A1 => net51553, A2 => net55953, ZN => net52292);
   U238 : NAND2_X1 port map( A1 => net51553, A2 => net55953, ZN => net47109);
   U239 : NAND2_X1 port map( A1 => DATA1(13), A2 => net46854, ZN => n306);
   U240 : NOR2_X1 port map( A1 => net55828, A2 => net46850, ZN => n308);
   U241 : AOI221_X1 port map( B1 => DATA1(6), B2 => n8, C1 => DATA1(14), C2 => 
                           net56098, A => n321, ZN => n323);
   U242 : INV_X1 port map( A => net50901, ZN => net50899);
   U243 : INV_X1 port map( A => DATA1(0), ZN => n139);
   U244 : INV_X1 port map( A => DATA1(16), ZN => n204);
   U245 : AOI22_X1 port map( A1 => n32, A2 => DATA1(8), B1 => net56281, B2 => 
                           DATA1(24), ZN => n49);
   U246 : NAND2_X1 port map( A1 => n113, A2 => net50839, ZN => n83);
   U247 : INV_X1 port map( A => n83, ZN => n50);
   U248 : NAND2_X1 port map( A1 => n50, A2 => net50869, ZN => n75);
   U249 : INV_X1 port map( A => n75, ZN => n51);
   U250 : NAND3_X1 port map( A1 => net50905, A2 => n51, A3 => net56256, ZN => 
                           n72);
   U251 : INV_X1 port map( A => DATA1(8), ZN => n258);
   U252 : OAI22_X1 port map( A1 => n258, A2 => net52292, B1 => n139, B2 => 
                           net56276, ZN => n52);
   U253 : INV_X1 port map( A => DATA1(4), ZN => n180);
   U254 : INV_X1 port map( A => DATA1(20), ZN => n298);
   U255 : AOI22_X1 port map( A1 => net55611, A2 => DATA1(12), B1 => n7, B2 => 
                           DATA1(28), ZN => n53);
   U256 : OAI221_X1 port map( B1 => net56277, B2 => n180, C1 => n298, C2 => 
                           net47197, A => n53, ZN => n76);
   U257 : INV_X1 port map( A => n76, ZN => n54);
   U258 : INV_X1 port map( A => DATA1(2), ZN => n161);
   U259 : INV_X1 port map( A => DATA1(10), ZN => n212);
   U260 : AOI22_X1 port map( A1 => net56281, A2 => DATA1(18), B1 => n7, B2 => 
                           DATA1(26), ZN => n56);
   U261 : OAI221_X1 port map( B1 => n161, B2 => net56277, C1 => n212, C2 => 
                           net52292, A => n56, ZN => n59);
   U262 : INV_X1 port map( A => DATA1(30), ZN => n320);
   U263 : NAND3_X1 port map( A1 => net55991, A2 => DATA1(6), A3 => net51553, ZN
                           => n58);
   U264 : AOI22_X1 port map( A1 => net56281, A2 => DATA1(22), B1 => net55611, 
                           B2 => DATA1(14), ZN => n57);
   U265 : OAI211_X1 port map( C1 => n320, C2 => n66, A => n58, B => n57, ZN => 
                           n93);
   U266 : MUX2_X1 port map( A => n59, B => n93, S => net50827, Z => n60);
   U267 : INV_X1 port map( A => n60, ZN => n78);
   U268 : INV_X1 port map( A => DATA1(9), ZN => n269);
   U269 : INV_X1 port map( A => DATA1(1), ZN => n150);
   U270 : OAI22_X1 port map( A1 => n269, A2 => net52292, B1 => n150, B2 => 
                           net47150, ZN => n62);
   U271 : INV_X1 port map( A => DATA1(5), ZN => net47043);
   U272 : INV_X1 port map( A => DATA1(29), ZN => net46850);
   U273 : NOR2_X1 port map( A1 => net56027, A2 => net46850, ZN => n63);
   U274 : AOI22_X1 port map( A1 => n63, A2 => net56120, B1 => net56225, B2 => 
                           DATA1(21), ZN => net47184);
   U275 : INV_X1 port map( A => net47157, ZN => net47183);
   U276 : MUX2_X1 port map( A => n64, B => net47183, S => net50827, Z => n69);
   U277 : AOI22_X1 port map( A1 => net56281, A2 => DATA1(19), B1 => n7, B2 => 
                           DATA1(27), ZN => n65);
   U278 : OAI221_X1 port map( B1 => net46879, B2 => net56277, C1 => net46973, 
                           C2 => net52292, A => n65, ZN => n67);
   U279 : OAI211_X1 port map( C1 => net46817, C2 => n66, A => net47177, B => 
                           net47178, ZN => n103);
   U280 : MUX2_X1 port map( A => n67, B => n103, S => net50827, Z => n68);
   U281 : INV_X1 port map( A => n68, ZN => n86);
   U282 : MUX2_X1 port map( A => n70, B => n79, S => net50889, Z => n71);
   U283 : NAND2_X1 port map( A1 => n72, A2 => n71, ZN => OUTPUT(0));
   U284 : INV_X1 port map( A => DATA1(17), ZN => n208);
   U285 : AOI22_X1 port map( A1 => n32, A2 => DATA1(9), B1 => net55672, B2 => 
                           DATA1(25), ZN => n73);
   U286 : OAI221_X1 port map( B1 => net55654, B2 => n150, C1 => n208, C2 => 
                           net47109, A => n73, ZN => n123);
   U287 : NAND2_X1 port map( A1 => n26, A2 => net50839, ZN => n91);
   U288 : INV_X1 port map( A => n91, ZN => n74);
   U289 : NAND2_X1 port map( A1 => n74, A2 => net50871, ZN => n84);
   U290 : MUX2_X1 port map( A => n84, B => n75, S => net50889, Z => n81);
   U291 : MUX2_X1 port map( A => n76, B => n113, S => net50827, Z => n77);
   U292 : INV_X1 port map( A => n77, ZN => n95);
   U293 : OAI22_X1 port map( A1 => net51547, A2 => n81, B1 => n80, B2 => 
                           net52168, ZN => OUTPUT(1));
   U294 : AOI22_X1 port map( A1 => net55611, A2 => DATA1(18), B1 => net56281, 
                           B2 => DATA1(26), ZN => n82);
   U295 : NAND2_X1 port map( A1 => n132, A2 => net50839, ZN => n101);
   U296 : MUX2_X1 port map( A => n101, B => n83, S => net50857, Z => n92);
   U297 : MUX2_X1 port map( A => n92, B => n84, S => net50889, Z => n89);
   U298 : INV_X1 port map( A => n85, ZN => n105);
   U299 : OAI22_X1 port map( A1 => net51553, A2 => n89, B1 => n88, B2 => 
                           net51543, ZN => OUTPUT(2));
   U300 : AOI22_X1 port map( A1 => n37, A2 => DATA1(19), B1 => net55672, B2 => 
                           DATA1(27), ZN => n90);
   U301 : OAI221_X1 port map( B1 => net55654, B2 => net46879, C1 => net46973, 
                           C2 => net56276, A => n90, ZN => n143);
   U302 : NAND2_X1 port map( A1 => n28, A2 => net50839, ZN => n111);
   U303 : MUX2_X1 port map( A => n111, B => n91, S => net50857, Z => n102);
   U304 : MUX2_X1 port map( A => n102, B => n92, S => net50889, Z => n98);
   U305 : MUX2_X1 port map( A => n93, B => n43, S => net50827, Z => n94);
   U306 : INV_X1 port map( A => n94, ZN => n115);
   U307 : MUX2_X1 port map( A => n95, B => n115, S => net50857, Z => n106);
   U308 : MUX2_X1 port map( A => n96, B => n106, S => net50889, Z => n97);
   U309 : OAI22_X1 port map( A1 => net51553, A2 => n98, B1 => n97, B2 => 
                           net51543, ZN => OUTPUT(3));
   U310 : AOI22_X1 port map( A1 => net56216, A2 => DATA1(12), B1 => net55672, 
                           B2 => DATA1(28), ZN => n99);
   U311 : OAI221_X1 port map( B1 => net55829, B2 => n180, C1 => n298, C2 => 
                           net52292, A => n99, ZN => n154);
   U312 : MUX2_X1 port map( A => n154, B => n113, S => net50827, Z => n100);
   U313 : INV_X1 port map( A => n100, ZN => n121);
   U314 : MUX2_X1 port map( A => n121, B => n101, S => net50857, Z => n112);
   U315 : MUX2_X1 port map( A => n112, B => n102, S => net50889, Z => n108);
   U316 : INV_X1 port map( A => n104, ZN => n125);
   U317 : OAI22_X1 port map( A1 => net51553, A2 => n108, B1 => n107, B2 => 
                           net51543, ZN => OUTPUT(4));
   U318 : INV_X1 port map( A => DATA1(21), ZN => net46851);
   U319 : AOI22_X1 port map( A1 => net56216, A2 => DATA1(13), B1 => net55672, 
                           B2 => DATA1(29), ZN => n109);
   U320 : OAI221_X1 port map( B1 => net55829, B2 => net47043, C1 => net46851, 
                           C2 => net47109, A => n109, ZN => n165);
   U321 : MUX2_X1 port map( A => n165, B => n123, S => net50827, Z => n110);
   U322 : INV_X1 port map( A => n110, ZN => n130);
   U323 : MUX2_X1 port map( A => n130, B => n111, S => net50857, Z => n122);
   U324 : MUX2_X1 port map( A => n122, B => n112, S => net50889, Z => n118);
   U325 : INV_X1 port map( A => n114, ZN => n134);
   U326 : MUX2_X1 port map( A => n116, B => n126, S => net50889, Z => n117);
   U327 : OAI22_X1 port map( A1 => net51551, A2 => n118, B1 => n117, B2 => 
                           net51543, ZN => OUTPUT(5));
   U328 : INV_X1 port map( A => DATA1(6), ZN => n194);
   U329 : INV_X1 port map( A => DATA1(22), ZN => n319);
   U330 : AOI22_X1 port map( A1 => n32, A2 => DATA1(14), B1 => net55672, B2 => 
                           DATA1(30), ZN => n119);
   U331 : OAI221_X1 port map( B1 => net55829, B2 => n194, C1 => n319, C2 => 
                           net47109, A => n119, ZN => n174);
   U332 : MUX2_X1 port map( A => n174, B => n132, S => net50827, Z => n120);
   U333 : INV_X1 port map( A => n120, ZN => n141);
   U334 : MUX2_X1 port map( A => n141, B => n121, S => net50857, Z => n131);
   U335 : MUX2_X1 port map( A => n131, B => n122, S => net50889, Z => n128);
   U336 : MUX2_X1 port map( A => n123, B => n165, S => net50833, Z => n124);
   U337 : INV_X1 port map( A => n124, ZN => n145);
   U338 : MUX2_X1 port map( A => n125, B => n145, S => net50857, Z => n135);
   U339 : OAI22_X1 port map( A1 => net51551, A2 => n128, B1 => n127, B2 => 
                           net51543, ZN => OUTPUT(6));
   U340 : MUX2_X1 port map( A => net47050, B => n143, S => net50831, Z => n129)
                           ;
   U341 : INV_X1 port map( A => n129, ZN => n152);
   U342 : MUX2_X1 port map( A => n152, B => n130, S => net50863, Z => n142);
   U343 : MUX2_X1 port map( A => n142, B => n131, S => net50891, Z => n137);
   U344 : MUX2_X1 port map( A => n43, B => n174, S => net50835, Z => n133);
   U345 : INV_X1 port map( A => n133, ZN => n156);
   U346 : MUX2_X1 port map( A => n135, B => n146, S => net50891, Z => n136);
   U347 : OAI22_X1 port map( A1 => net51551, A2 => n137, B1 => n136, B2 => 
                           net51543, ZN => OUTPUT(7));
   U348 : AOI22_X1 port map( A1 => net55611, A2 => DATA1(24), B1 => net56216, 
                           B2 => DATA1(16), ZN => n138);
   U349 : MUX2_X1 port map( A => net47039, B => n154, S => net50833, Z => n140)
                           ;
   U350 : INV_X1 port map( A => n140, ZN => n163);
   U351 : MUX2_X1 port map( A => n163, B => n141, S => net50857, Z => n153);
   U352 : MUX2_X1 port map( A => n153, B => n142, S => net50891, Z => n148);
   U353 : MUX2_X1 port map( A => n143, B => net47050, S => net50835, Z => n144)
                           ;
   U354 : INV_X1 port map( A => n144, ZN => n167);
   U355 : OAI22_X1 port map( A1 => net51551, A2 => n148, B1 => n147, B2 => 
                           net51543, ZN => OUTPUT(8));
   U356 : AOI22_X1 port map( A1 => n37, A2 => DATA1(25), B1 => DATA1(17), B2 =>
                           n32, ZN => n149);
   U357 : OAI221_X1 port map( B1 => n150, B2 => net51703, C1 => net51599, C2 =>
                           n269, A => n149, ZN => net47028);
   U358 : MUX2_X1 port map( A => net47028, B => n165, S => n9, Z => n151);
   U359 : INV_X1 port map( A => n151, ZN => n172);
   U360 : MUX2_X1 port map( A => n172, B => n152, S => net50861, Z => n164);
   U361 : MUX2_X1 port map( A => n164, B => n153, S => net50891, Z => n159);
   U362 : MUX2_X1 port map( A => n154, B => n46, S => n9, Z => n155);
   U363 : INV_X1 port map( A => n155, ZN => n175);
   U364 : MUX2_X1 port map( A => n157, B => n168, S => net50891, Z => n158);
   U365 : OAI22_X1 port map( A1 => net51551, A2 => n159, B1 => n158, B2 => 
                           net51543, ZN => OUTPUT(9));
   U366 : AOI22_X1 port map( A1 => n37, A2 => DATA1(26), B1 => n32, B2 => 
                           DATA1(18), ZN => n160);
   U367 : OAI221_X1 port map( B1 => net55829, B2 => n212, C1 => net56284, C2 =>
                           n161, A => n160, ZN => n201);
   U368 : MUX2_X1 port map( A => n201, B => n174, S => net50833, Z => n162);
   U369 : INV_X1 port map( A => n162, ZN => n182);
   U370 : MUX2_X1 port map( A => n182, B => n163, S => net50865, Z => n173);
   U371 : MUX2_X1 port map( A => n173, B => n164, S => net50891, Z => n170);
   U372 : MUX2_X1 port map( A => n165, B => net47028, S => n9, Z => n166);
   U373 : INV_X1 port map( A => n166, ZN => n184);
   U374 : MUX2_X1 port map( A => n167, B => n184, S => net50857, Z => n176);
   U375 : OAI22_X1 port map( A1 => net51551, A2 => n170, B1 => n169, B2 => 
                           net51543, ZN => OUTPUT(10));
   U376 : AOI22_X1 port map( A1 => n37, A2 => DATA1(27), B1 => net56178, B2 => 
                           DATA1(19), ZN => net47065);
   U377 : MUX2_X1 port map( A => net56186, B => net47050, S => net50831, Z => 
                           n171);
   U378 : INV_X1 port map( A => n171, ZN => n188);
   U379 : MUX2_X1 port map( A => n188, B => n172, S => net50857, Z => n183);
   U380 : MUX2_X1 port map( A => n183, B => n173, S => net50891, Z => n178);
   U381 : MUX2_X1 port map( A => n174, B => n201, S => net50835, Z => net47060)
                           ;
   U382 : INV_X1 port map( A => net47060, ZN => net47037);
   U383 : MUX2_X1 port map( A => n176, B => n185, S => net50891, Z => n177);
   U384 : OAI22_X1 port map( A1 => net51551, A2 => n178, B1 => n177, B2 => 
                           net51543, ZN => OUTPUT(11));
   U385 : INV_X1 port map( A => DATA1(12), ZN => n223);
   U386 : AOI22_X1 port map( A1 => n37, A2 => DATA1(28), B1 => n32, B2 => 
                           DATA1(20), ZN => n179);
   U387 : OAI221_X1 port map( B1 => net56146, B2 => n180, C1 => net56118, C2 =>
                           n223, A => n179, ZN => n209);
   U388 : MUX2_X1 port map( A => n209, B => n46, S => net50835, Z => n181);
   U389 : INV_X1 port map( A => n181, ZN => n196);
   U390 : MUX2_X1 port map( A => n196, B => n182, S => net50865, Z => n189);
   U391 : MUX2_X1 port map( A => n189, B => n183, S => net50891, Z => n187);
   U392 : INV_X1 port map( A => net47049, ZN => net47026);
   U393 : OAI22_X1 port map( A1 => net51549, A2 => n187, B1 => n186, B2 => 
                           net51543, ZN => OUTPUT(12));
   U394 : INV_X1 port map( A => net47042, ZN => net47018);
   U395 : MUX2_X1 port map( A => net47018, B => n188, S => net50861, Z => n197)
                           ;
   U396 : MUX2_X1 port map( A => n197, B => n189, S => net50893, Z => n192);
   U397 : OAI22_X1 port map( A1 => net51549, A2 => n192, B1 => n191, B2 => 
                           net51543, ZN => OUTPUT(13));
   U398 : INV_X1 port map( A => DATA1(14), ZN => n240);
   U399 : AOI22_X1 port map( A1 => net55611, A2 => DATA1(30), B1 => net56216, 
                           B2 => DATA1(22), ZN => n193);
   U400 : MUX2_X1 port map( A => net56195, B => net56192, S => net50831, Z => 
                           n195);
   U401 : INV_X1 port map( A => n195, ZN => n206);
   U402 : MUX2_X1 port map( A => n206, B => n196, S => net50861, Z => n200);
   U403 : MUX2_X1 port map( A => n200, B => n197, S => net50893, Z => n199);
   U404 : OAI22_X1 port map( A1 => net51549, A2 => n199, B1 => n198, B2 => 
                           net51543, ZN => OUTPUT(14));
   U405 : INV_X1 port map( A => net47019, ZN => net46994);
   U406 : MUX2_X1 port map( A => net46994, B => net47018, S => net50861, Z => 
                           net47004);
   U407 : MUX2_X1 port map( A => net47004, B => n200, S => net50893, Z => n202)
                           ;
   U408 : OAI22_X1 port map( A1 => net51549, A2 => n202, B1 => net47012, B2 => 
                           net51543, ZN => OUTPUT(15));
   U409 : NAND2_X1 port map( A1 => net55782, A2 => net55980, ZN => net47009);
   U410 : INV_X1 port map( A => net47009, ZN => net46854);
   U411 : AOI22_X1 port map( A1 => n12, A2 => DATA1(0), B1 => net56216, B2 => 
                           DATA1(24), ZN => n203);
   U412 : OAI221_X1 port map( B1 => n258, B2 => net51703, C1 => net56118, C2 =>
                           n204, A => n203, ZN => n233);
   U413 : MUX2_X1 port map( A => n233, B => net55789, S => net50831, Z => n205)
                           ;
   U414 : INV_X1 port map( A => n205, ZN => n214);
   U415 : AOI22_X1 port map( A1 => n11, A2 => DATA1(1), B1 => net56216, B2 => 
                           DATA1(25), ZN => n207);
   U416 : OAI221_X1 port map( B1 => n10, B2 => n269, C1 => net56118, C2 => n208
                           , A => n207, ZN => net46936);
   U417 : INV_X1 port map( A => net46995, ZN => net46971);
   U418 : MUX2_X1 port map( A => net46971, B => net46994, S => net50861, Z => 
                           n215);
   U419 : MUX2_X1 port map( A => n215, B => net46993, S => net50893, Z => n210)
                           ;
   U420 : MUX2_X1 port map( A => n209, B => n233, S => net50831, Z => net46991)
                           ;
   U421 : INV_X1 port map( A => net46991, ZN => net46967);
   U422 : OAI22_X1 port map( A1 => net51549, A2 => n210, B1 => net46988, B2 => 
                           net51543, ZN => OUTPUT(17));
   U423 : INV_X1 port map( A => DATA1(18), ZN => n280);
   U424 : AOI22_X1 port map( A1 => n11, A2 => DATA1(2), B1 => net56216, B2 => 
                           DATA1(26), ZN => n211);
   U425 : MUX2_X1 port map( A => n33, B => net56195, S => net50831, Z => n213);
   U426 : INV_X1 port map( A => n213, ZN => n225);
   U427 : MUX2_X1 port map( A => n225, B => n214, S => net50861, Z => n218);
   U428 : MUX2_X1 port map( A => n218, B => n215, S => net50893, Z => n217);
   U429 : INV_X1 port map( A => net46980, ZN => net46956);
   U430 : OAI22_X1 port map( A1 => net51547, A2 => n217, B1 => n216, B2 => 
                           net51543, ZN => OUTPUT(18));
   U431 : INV_X1 port map( A => DATA1(19), ZN => net46974);
   U432 : OAI221_X1 port map( B1 => n10, B2 => net46973, C1 => net51599, C2 => 
                           net46974, A => net46975, ZN => net46911);
   U433 : INV_X1 port map( A => net46972, ZN => net46949);
   U434 : MUX2_X1 port map( A => net46949, B => net46971, S => net50863, Z => 
                           n226);
   U435 : MUX2_X1 port map( A => n226, B => n218, S => net50895, Z => n221);
   U436 : INV_X1 port map( A => n219, ZN => n235);
   U437 : MUX2_X1 port map( A => net46966, B => n227, S => net50895, Z => n220)
                           ;
   U438 : OAI22_X1 port map( A1 => net51547, A2 => n221, B1 => n220, B2 => 
                           net51543, ZN => OUTPUT(19));
   U439 : AOI22_X1 port map( A1 => DATA1(4), A2 => net55740, B1 => net56178, B2
                           => DATA1(28), ZN => n222);
   U440 : OAI221_X1 port map( B1 => n10, B2 => n223, C1 => net51599, C2 => n298
                           , A => n222, ZN => n273);
   U441 : MUX2_X1 port map( A => n273, B => n233, S => net50833, Z => n224);
   U442 : INV_X1 port map( A => n224, ZN => n242);
   U443 : MUX2_X1 port map( A => n242, B => n225, S => net50863, Z => n232);
   U444 : MUX2_X1 port map( A => n232, B => n226, S => net50895, Z => n229);
   U445 : INV_X1 port map( A => net46957, ZN => net46934);
   U446 : OAI22_X1 port map( A1 => net51547, A2 => n229, B1 => n228, B2 => 
                           net56256, ZN => OUTPUT(20));
   U447 : AOI22_X1 port map( A1 => DATA1(5), A2 => net55741, B1 => net56178, B2
                           => DATA1(29), ZN => n230);
   U448 : MUX2_X1 port map( A => n30, B => net46936, S => net50833, Z => n231);
   U449 : INV_X1 port map( A => n231, ZN => n249);
   U450 : MUX2_X1 port map( A => n249, B => net46949, S => net50863, Z => n243)
                           ;
   U451 : MUX2_X1 port map( A => n243, B => n232, S => net50895, Z => n238);
   U452 : INV_X1 port map( A => n234, ZN => n252);
   U453 : OAI22_X1 port map( A1 => net51547, A2 => n238, B1 => n237, B2 => 
                           net56256, ZN => OUTPUT(21));
   U454 : AOI22_X1 port map( A1 => net55739, A2 => DATA1(6), B1 => net56178, B2
                           => DATA1(30), ZN => n239);
   U455 : OAI221_X1 port map( B1 => n10, B2 => n240, C1 => net55828, C2 => n319
                           , A => n239, ZN => n291);
   U456 : MUX2_X1 port map( A => n291, B => n33, S => net50833, Z => n241);
   U457 : INV_X1 port map( A => n241, ZN => n260);
   U458 : MUX2_X1 port map( A => n260, B => n242, S => net50863, Z => n250);
   U459 : MUX2_X1 port map( A => n250, B => n243, S => net50895, Z => n247);
   U460 : INV_X1 port map( A => n244, ZN => n263);
   U461 : OAI22_X1 port map( A1 => net51547, A2 => n247, B1 => n246, B2 => 
                           net56256, ZN => OUTPUT(22));
   U462 : MUX2_X1 port map( A => net46859, B => net46911, S => net50833, Z => 
                           n248);
   U463 : INV_X1 port map( A => n248, ZN => n271);
   U464 : MUX2_X1 port map( A => n261, B => n250, S => net50895, Z => n255);
   U465 : INV_X1 port map( A => n251, ZN => n274);
   U466 : OAI22_X1 port map( A1 => net51549, A2 => n255, B1 => n254, B2 => 
                           net52168, ZN => OUTPUT(23));
   U467 : NAND3_X1 port map( A1 => DATA1(24), A2 => net55100, A3 => net52169, 
                           ZN => n257);
   U468 : AOI22_X1 port map( A1 => DATA1(16), A2 => net46881, B1 => DATA1(0), 
                           B2 => n8, ZN => n256);
   U469 : OAI211_X1 port map( C1 => net46901, C2 => n258, A => n257, B => n256,
                           ZN => n299);
   U470 : MUX2_X1 port map( A => n299, B => n273, S => net50833, Z => n259);
   U471 : INV_X1 port map( A => n259, ZN => n282);
   U472 : MUX2_X1 port map( A => n282, B => n260, S => net50863, Z => n272);
   U473 : MUX2_X1 port map( A => n272, B => n261, S => net50895, Z => n266);
   U474 : INV_X1 port map( A => n262, ZN => n284);
   U475 : OAI22_X1 port map( A1 => net51547, A2 => n266, B1 => n265, B2 => 
                           net51543, ZN => OUTPUT(24));
   U476 : NAND3_X1 port map( A1 => DATA1(25), A2 => net55991, A3 => net52169, 
                           ZN => n268);
   U477 : AOI22_X1 port map( A1 => DATA1(17), A2 => net46881, B1 => DATA1(1), 
                           B2 => n8, ZN => n267);
   U478 : MUX2_X1 port map( A => n29, B => n30, S => net50835, Z => n270);
   U479 : INV_X1 port map( A => n270, ZN => n289);
   U480 : MUX2_X1 port map( A => n289, B => n271, S => net50865, Z => n283);
   U481 : MUX2_X1 port map( A => n283, B => n272, S => net50897, Z => n277);
   U482 : NAND2_X1 port map( A1 => n273, A2 => net50839, ZN => n292);
   U483 : MUX2_X1 port map( A => n275, B => n285, S => net50897, Z => n276);
   U484 : OAI22_X1 port map( A1 => net51547, A2 => n277, B1 => n276, B2 => 
                           net56256, ZN => OUTPUT(25));
   U485 : INV_X1 port map( A => DATA1(26), ZN => n279);
   U486 : AOI22_X1 port map( A1 => DATA1(10), A2 => net55739, B1 => DATA1(2), 
                           B2 => n8, ZN => n278);
   U487 : MUX2_X1 port map( A => n322, B => n291, S => net50835, Z => n281);
   U488 : INV_X1 port map( A => n281, ZN => n302);
   U489 : MUX2_X1 port map( A => n302, B => n282, S => net50865, Z => n290);
   U490 : MUX2_X1 port map( A => n290, B => n283, S => net50897, Z => n287);
   U491 : NAND2_X1 port map( A1 => n30, A2 => net50841, ZN => n304);
   U492 : MUX2_X1 port map( A => n284, B => n304, S => net50865, Z => n293);
   U493 : OAI22_X1 port map( A1 => net51549, A2 => n287, B1 => n286, B2 => 
                           net56256, ZN => OUTPUT(26));
   U494 : INV_X1 port map( A => DATA1(27), ZN => net46877);
   U495 : OAI221_X1 port map( B1 => net55828, B2 => net46877, C1 => net46878, 
                           C2 => net46879, A => net46880, ZN => n331);
   U496 : MUX2_X1 port map( A => n331, B => net46859, S => net50835, Z => n288)
                           ;
   U497 : INV_X1 port map( A => n288, ZN => n313);
   U498 : MUX2_X1 port map( A => n303, B => n290, S => net50897, Z => n295);
   U499 : NAND2_X1 port map( A1 => n36, A2 => net50841, ZN => n315);
   U500 : MUX2_X1 port map( A => n292, B => n315, S => net50865, Z => net46857)
                           ;
   U501 : MUX2_X1 port map( A => n293, B => net46857, S => net50897, Z => n294)
                           ;
   U502 : OAI22_X1 port map( A1 => net51549, A2 => n295, B1 => n294, B2 => 
                           net56256, ZN => OUTPUT(27));
   U503 : INV_X1 port map( A => DATA1(28), ZN => n297);
   U504 : AOI22_X1 port map( A1 => DATA1(4), A2 => n8, B1 => net55741, B2 => 
                           DATA1(12), ZN => n296);
   U505 : MUX2_X1 port map( A => n300, B => n299, S => net50835, Z => n301);
   U506 : INV_X1 port map( A => n301, ZN => n324);
   U507 : MUX2_X1 port map( A => n324, B => n302, S => net50865, Z => n314);
   U508 : MUX2_X1 port map( A => n314, B => n303, S => net50897, Z => n305);
   U509 : NAND2_X1 port map( A1 => net55902, A2 => net50841, ZN => n327);
   U510 : OAI22_X1 port map( A1 => n305, A2 => net51551, B1 => net46856, B2 => 
                           net56256, ZN => OUTPUT(28));
   U511 : NAND3_X1 port map( A1 => DATA1(5), A2 => n1, A3 => net56120, ZN => 
                           n307);
   U512 : MUX2_X1 port map( A => n333, B => n313, S => net50865, Z => n326);
   U513 : MUX2_X1 port map( A => n35, B => n314, S => net50897, Z => n318);
   U514 : INV_X1 port map( A => n315, ZN => n316);
   U515 : NAND2_X1 port map( A1 => n316, A2 => net50871, ZN => n328);
   U516 : MUX2_X1 port map( A => net46838, B => n328, S => net50897, Z => n317)
                           ;
   U517 : OAI22_X1 port map( A1 => n318, A2 => net51549, B1 => n317, B2 => 
                           net52168, ZN => OUTPUT(29));
   U518 : OAI22_X1 port map( A1 => net55828, A2 => n320, B1 => n319, B2 => 
                           net51702, ZN => n321);
   U519 : MUX2_X1 port map( A => n325, B => n324, S => net50865, Z => n335);
   U520 : NAND2_X1 port map( A1 => n3, A2 => net50871, ZN => n337);
   U521 : MUX2_X1 port map( A => n328, B => n337, S => net50899, Z => n329);
   U522 : OAI22_X1 port map( A1 => n330, A2 => net51549, B1 => n329, B2 => 
                           net52168, ZN => OUTPUT(30));
   U523 : OAI22_X1 port map( A1 => net55828, A2 => net46817, B1 => net51702, B2
                           => net46819, ZN => net46815);
   U524 : INV_X1 port map( A => n331, ZN => n332);
   U525 : MUX2_X1 port map( A => net46810, B => n332, S => net50835, Z => n334)
                           ;
   U526 : MUX2_X1 port map( A => n334, B => n333, S => net50865, Z => n336);
   U527 : MUX2_X1 port map( A => n336, B => n335, S => net50899, Z => n340);
   U528 : INV_X1 port map( A => n337, ZN => n338);
   U529 : NAND3_X1 port map( A1 => net50905, A2 => n338, A3 => net51553, ZN => 
                           n339);
   U530 : NAND2_X1 port map( A1 => n340, A2 => n339, ZN => OUTPUT(31));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_0 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_0;

architecture SYN_BEHAVIOUR of NAND4_0 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => B, A2 => A, A3 => D, A4 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_96 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_96;

architecture SYN_BEHAVIOUR of NAND3_96 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_0 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_0;

architecture SYN_BEHAVIOUR of NAND3_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_N32_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end ADDER_N32_DW01_add_0;

architecture SYN_rpl of ADDER_N32_DW01_add_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port, 
      SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, SUM_17_port, 
      SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, 
      SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, SUM_30_port, SUM_31_port, SUM_3_port, 
      SUM_4_port, SUM_5_port, SUM_6_port, SUM_7_port, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : XOR2_X1 port map( A => A(8), B => n34, Z => SUM_8_port);
   U2 : XOR2_X1 port map( A => A(9), B => n35, Z => SUM_9_port);
   U3 : XOR2_X1 port map( A => A(10), B => n36, Z => SUM_10_port);
   U4 : XOR2_X1 port map( A => A(11), B => n37, Z => SUM_11_port);
   U5 : XOR2_X1 port map( A => A(12), B => n38, Z => SUM_12_port);
   U6 : XOR2_X1 port map( A => A(13), B => n39, Z => SUM_13_port);
   U7 : XOR2_X1 port map( A => A(14), B => n40, Z => SUM_14_port);
   U8 : XOR2_X1 port map( A => A(15), B => n41, Z => SUM_15_port);
   U9 : XOR2_X1 port map( A => A(16), B => n42, Z => SUM_16_port);
   U10 : XOR2_X1 port map( A => A(17), B => n43, Z => SUM_17_port);
   U11 : XOR2_X1 port map( A => A(18), B => n44, Z => SUM_18_port);
   U12 : XOR2_X1 port map( A => A(19), B => n45, Z => SUM_19_port);
   U13 : XOR2_X1 port map( A => A(20), B => n46, Z => SUM_20_port);
   U14 : XOR2_X1 port map( A => A(21), B => n47, Z => SUM_21_port);
   U15 : XOR2_X1 port map( A => A(22), B => n48, Z => SUM_22_port);
   U16 : XOR2_X1 port map( A => A(23), B => n49, Z => SUM_23_port);
   U17 : XOR2_X1 port map( A => A(24), B => n50, Z => SUM_24_port);
   U18 : XOR2_X1 port map( A => A(25), B => n51, Z => SUM_25_port);
   U19 : XOR2_X1 port map( A => A(26), B => n52, Z => SUM_26_port);
   U20 : XOR2_X1 port map( A => A(27), B => n53, Z => SUM_27_port);
   U21 : XOR2_X1 port map( A => A(28), B => n54, Z => SUM_28_port);
   U22 : XOR2_X1 port map( A => A(29), B => n55, Z => SUM_29_port);
   U23 : XOR2_X1 port map( A => A(30), B => n56, Z => SUM_30_port);
   U24 : XOR2_X1 port map( A => A(31), B => n57, Z => SUM_31_port);
   U25 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U26 : XOR2_X1 port map( A => A(4), B => n30, Z => SUM_4_port);
   U27 : XOR2_X1 port map( A => A(5), B => n31, Z => SUM_5_port);
   U28 : XOR2_X1 port map( A => A(6), B => n32, Z => SUM_6_port);
   U29 : XOR2_X1 port map( A => A(7), B => n33, Z => SUM_7_port);
   U30 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n30);
   U31 : AND2_X1 port map( A1 => A(4), A2 => n30, ZN => n31);
   U32 : AND2_X1 port map( A1 => A(5), A2 => n31, ZN => n32);
   U33 : AND2_X1 port map( A1 => A(6), A2 => n32, ZN => n33);
   U34 : AND2_X1 port map( A1 => A(7), A2 => n33, ZN => n34);
   U35 : AND2_X1 port map( A1 => A(8), A2 => n34, ZN => n35);
   U36 : AND2_X1 port map( A1 => A(9), A2 => n35, ZN => n36);
   U37 : AND2_X1 port map( A1 => A(10), A2 => n36, ZN => n37);
   U38 : AND2_X1 port map( A1 => A(11), A2 => n37, ZN => n38);
   U39 : AND2_X1 port map( A1 => A(12), A2 => n38, ZN => n39);
   U40 : AND2_X1 port map( A1 => A(13), A2 => n39, ZN => n40);
   U41 : AND2_X1 port map( A1 => A(14), A2 => n40, ZN => n41);
   U42 : AND2_X1 port map( A1 => A(15), A2 => n41, ZN => n42);
   U43 : AND2_X1 port map( A1 => A(16), A2 => n42, ZN => n43);
   U44 : AND2_X1 port map( A1 => A(17), A2 => n43, ZN => n44);
   U45 : AND2_X1 port map( A1 => A(18), A2 => n44, ZN => n45);
   U46 : AND2_X1 port map( A1 => A(19), A2 => n45, ZN => n46);
   U47 : AND2_X1 port map( A1 => A(20), A2 => n46, ZN => n47);
   U48 : AND2_X1 port map( A1 => A(21), A2 => n47, ZN => n48);
   U49 : AND2_X1 port map( A1 => A(22), A2 => n48, ZN => n49);
   U50 : AND2_X1 port map( A1 => A(23), A2 => n49, ZN => n50);
   U51 : AND2_X1 port map( A1 => A(24), A2 => n50, ZN => n51);
   U52 : AND2_X1 port map( A1 => A(25), A2 => n51, ZN => n52);
   U53 : AND2_X1 port map( A1 => A(26), A2 => n52, ZN => n53);
   U54 : AND2_X1 port map( A1 => A(27), A2 => n53, ZN => n54);
   U55 : AND2_X1 port map( A1 => A(28), A2 => n54, ZN => n55);
   U56 : AND2_X1 port map( A1 => A(29), A2 => n55, ZN => n56);
   U57 : AND2_X1 port map( A1 => A(30), A2 => n56, ZN => n57);
   U58 : INV_X1 port map( A => A(2), ZN => SUM_2_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32 is

   port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
         downto 0));

end ALU_N32;

architecture SYN_BEHAVIOR of ALU_N32 is

   component ALU_N32_DW01_cmp6_3
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component ALU_N32_DW01_cmp6_2
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component ALU_N32_DW01_add_2
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component ALU_N32_DW01_sub_2
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component BARREL_SHIFTER_N32
      port( CONF : in std_logic;  DATA1, DATA2 : in std_logic_vector (31 downto
            0);  OUTPUT : out std_logic_vector (31 downto 0));
   end component;
   
   component NAND4_1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_2
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_3
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_4
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_5
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_6
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_7
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_8
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_9
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_10
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_11
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_12
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_13
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_14
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_15
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_16
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_17
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_18
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_19
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_20
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_21
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_22
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_23
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_24
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_25
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_26
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_27
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_28
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_29
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_30
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_31
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_0
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_2
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_3
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_4
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_5
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_6
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_7
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_8
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_9
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_10
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_11
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_12
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_13
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_14
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_15
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_16
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_17
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_18
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_19
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_20
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_21
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_22
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_23
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_24
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_25
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_26
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_27
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_28
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_29
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_30
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_31
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_32
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_33
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_34
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_35
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_36
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_37
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_38
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_39
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_40
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_41
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_42
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_43
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_44
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_45
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_46
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_47
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_48
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_49
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_50
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_51
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_52
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_53
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_54
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_55
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_56
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_57
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_58
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_59
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_60
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_61
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_62
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_63
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_64
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_65
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_66
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_67
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_68
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_69
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_70
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_71
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_72
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_73
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_74
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_75
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_76
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_77
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_78
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_79
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_80
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_81
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_82
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_83
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_84
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_85
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_86
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_87
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_88
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_89
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_90
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_91
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_92
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_93
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_94
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_95
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_96
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_97
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_98
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_99
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_100
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_101
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_102
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_103
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_104
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_105
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_106
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_107
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_108
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_109
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_110
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_111
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_112
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_113
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_114
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_115
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_116
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_117
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_118
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_119
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_120
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_121
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_122
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_123
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_124
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_125
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_126
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_127
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_0
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
      N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72
      , N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, 
      N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, 
      N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, 
      Y_LOGIC_31_port, Y_LOGIC_30_port, Y_LOGIC_29_port, Y_LOGIC_28_port, 
      Y_LOGIC_27_port, Y_LOGIC_26_port, Y_LOGIC_25_port, Y_LOGIC_24_port, 
      Y_LOGIC_23_port, Y_LOGIC_22_port, Y_LOGIC_21_port, Y_LOGIC_20_port, 
      Y_LOGIC_19_port, Y_LOGIC_18_port, Y_LOGIC_17_port, Y_LOGIC_16_port, 
      Y_LOGIC_15_port, Y_LOGIC_14_port, Y_LOGIC_13_port, Y_LOGIC_12_port, 
      Y_LOGIC_11_port, Y_LOGIC_10_port, Y_LOGIC_9_port, Y_LOGIC_8_port, 
      Y_LOGIC_7_port, Y_LOGIC_6_port, Y_LOGIC_5_port, Y_LOGIC_4_port, 
      Y_LOGIC_3_port, Y_LOGIC_2_port, Y_LOGIC_1_port, Y_LOGIC_0_port, N111, 
      N112, N113, OUT_SHIFTER_31_port, OUT_SHIFTER_30_port, OUT_SHIFTER_29_port
      , OUT_SHIFTER_28_port, OUT_SHIFTER_27_port, OUT_SHIFTER_26_port, 
      OUT_SHIFTER_25_port, OUT_SHIFTER_24_port, OUT_SHIFTER_23_port, 
      OUT_SHIFTER_22_port, OUT_SHIFTER_21_port, OUT_SHIFTER_20_port, 
      OUT_SHIFTER_19_port, OUT_SHIFTER_18_port, OUT_SHIFTER_17_port, 
      OUT_SHIFTER_16_port, OUT_SHIFTER_15_port, OUT_SHIFTER_14_port, 
      OUT_SHIFTER_13_port, OUT_SHIFTER_12_port, OUT_SHIFTER_11_port, 
      OUT_SHIFTER_10_port, OUT_SHIFTER_9_port, OUT_SHIFTER_8_port, 
      OUT_SHIFTER_7_port, OUT_SHIFTER_6_port, OUT_SHIFTER_5_port, 
      OUT_SHIFTER_4_port, OUT_SHIFTER_3_port, OUT_SHIFTER_2_port, 
      OUT_SHIFTER_1_port, OUT_SHIFTER_0_port, S_3_port, L0_31_port, L0_30_port,
      L0_29_port, L0_28_port, L0_27_port, L0_26_port, L0_25_port, L0_24_port, 
      L0_23_port, L0_22_port, L0_21_port, L0_20_port, L0_19_port, L0_18_port, 
      L0_17_port, L0_16_port, L0_15_port, L0_14_port, L0_13_port, L0_12_port, 
      L0_11_port, L0_10_port, L0_9_port, L0_8_port, L0_7_port, L0_6_port, 
      L0_5_port, L0_4_port, L0_3_port, L0_2_port, L0_1_port, L0_0_port, 
      L1_31_port, L1_30_port, L1_29_port, L1_28_port, L1_27_port, L1_26_port, 
      L1_25_port, L1_24_port, L1_23_port, L1_22_port, L1_21_port, L1_20_port, 
      L1_19_port, L1_18_port, L1_17_port, L1_16_port, L1_15_port, L1_14_port, 
      L1_13_port, L1_12_port, L1_11_port, L1_10_port, L1_9_port, L1_8_port, 
      L1_7_port, L1_6_port, L1_5_port, L1_4_port, L1_3_port, L1_2_port, 
      L1_1_port, L1_0_port, L2_31_port, L2_30_port, L2_29_port, L2_28_port, 
      L2_27_port, L2_26_port, L2_25_port, L2_24_port, L2_23_port, L2_22_port, 
      L2_21_port, L2_20_port, L2_19_port, L2_18_port, L2_17_port, L2_16_port, 
      L2_15_port, L2_14_port, L2_13_port, L2_12_port, L2_11_port, L2_10_port, 
      L2_9_port, L2_8_port, L2_7_port, L2_6_port, L2_5_port, L2_4_port, 
      L2_3_port, L2_2_port, L2_1_port, L2_0_port, L3_31_port, L3_30_port, 
      L3_29_port, L3_28_port, L3_27_port, L3_26_port, L3_25_port, L3_24_port, 
      L3_23_port, L3_22_port, L3_21_port, L3_20_port, L3_19_port, L3_18_port, 
      L3_17_port, L3_16_port, L3_15_port, L3_14_port, L3_13_port, L3_12_port, 
      L3_11_port, L3_10_port, L3_9_port, L3_8_port, L3_7_port, L3_6_port, 
      L3_5_port, L3_4_port, L3_3_port, L3_2_port, L3_1_port, L3_0_port, n10, 
      n11, n12, n13, net23929, net47281, net47283, net47284, net47289, net47290
      , net47291, net51571, net51569, net51567, net51565, net51563, net51561, 
      net51577, net51575, net51573, net51583, net51581, net51579, net51589, 
      net51587, net51585, net51595, net51593, net51591, net51772, net54989, 
      net55526, net55932, net56011, net54984, net47243, net56205, net56055, 
      net55940, net47294, net47292, net47288, net47282, net47280, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47_port, n48_port, n49_port, 
      n50_port, n51_port, n52_port, n53_port, n54_port, n55_port, n56_port, 
      n57_port, n58_port, n59_port, n60_port, n61_port, n62_port, n63_port, 
      n64_port, n65_port, n66_port, n67_port, n68_port, n69_port, n70_port, 
      n71_port, n72_port, n73_port, n74_port, n75_port, n76_port, n77_port, 
      n78_port, n79_port, n80_port, n81_port, n82_port, n83_port, n84_port, 
      n85_port, n86_port, n87_port, n88_port, n89_port, n90_port, n91_port, 
      n92_port, n93_port, n94_port, n95_port, n96_port, n97_port, n98_port, 
      n99_port, n100_port, n101_port, n102_port, n103_port, n104_port, 
      n105_port, n106_port, n107_port, n108_port, n109_port, n110_port, 
      n111_port, n112_port, n113_port, n114, n115, n116, n117, n118, n119, n120
      , n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n_1150, n_1151, n_1152, n_1153,
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160 : std_logic;

begin
   
   X_Logic0_port <= '0';
   n10 <= '0';
   n11 <= '0';
   n12 <= '0';
   n13 <= '1';
   U5 : INV_X1 port map( A => n226, ZN => n1);
   U6 : CLKBUF_X1 port map( A => DATA1(1), Z => n129);
   U7 : BUF_X1 port map( A => net54984, Z => net51579);
   U8 : BUF_X1 port map( A => n18, Z => net51589);
   U10 : BUF_X1 port map( A => n21, Z => n32);
   U11 : BUF_X2 port map( A => n72_port, Z => n97_port);
   U12 : CLKBUF_X1 port map( A => FUNC(2), Z => n17);
   U13 : AND4_X2 port map( A1 => net56055, A2 => net47288, A3 => FUNC(0), A4 =>
                           FUNC(3), ZN => net55526);
   U14 : NAND2_X1 port map( A1 => N75, A2 => net51573, ZN => n2);
   U15 : AND2_X1 port map( A1 => Y_LOGIC_28_port, A2 => net51585, ZN => n4);
   U16 : NAND2_X1 port map( A1 => N107, A2 => net51579, ZN => n5);
   U17 : AND2_X1 port map( A1 => n5, A2 => n6, ZN => n3);
   U18 : AND2_X1 port map( A1 => n7, A2 => n2, ZN => n6);
   U19 : INV_X1 port map( A => n4, ZN => n7);
   U20 : NAND2_X1 port map( A1 => OUT_SHIFTER_16_port, A2 => net51593, ZN => n9
                           );
   U21 : NAND2_X1 port map( A1 => n9, A2 => net47243, ZN => OUTALU(16));
   U22 : BUF_X2 port map( A => n8, Z => net51593);
   U23 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n8);
   U24 : BUF_X2 port map( A => n8, Z => net51591);
   U25 : CLKBUF_X3 port map( A => n8, Z => net51595);
   U26 : NAND4_X1 port map( A1 => net56205, A2 => net55932, A3 => net55940, A4 
                           => net51772, ZN => n15);
   U27 : INV_X1 port map( A => n17, ZN => net51772);
   U28 : CLKBUF_X1 port map( A => n17, Z => n16);
   U29 : NAND3_X1 port map( A1 => n17, A2 => net55932, A3 => net54989, ZN => 
                           net47284);
   U30 : CLKBUF_X1 port map( A => net47292, Z => net55940);
   U31 : INV_X1 port map( A => net55940, ZN => net56011);
   U32 : OAI33_X1 port map( A1 => net47291, A2 => net55932, A3 => net47282, B1 
                           => net56205, B2 => net51772, B3 => net55940, ZN => 
                           net47290);
   U33 : INV_X1 port map( A => FUNC(1), ZN => net47292);
   U34 : AND2_X1 port map( A1 => net47294, A2 => net47292, ZN => net54989);
   U35 : NAND2_X1 port map( A1 => net56205, A2 => net47292, ZN => net47282);
   U36 : INV_X1 port map( A => net47281, ZN => net55932);
   U37 : INV_X1 port map( A => FUNC(3), ZN => net47281);
   U38 : INV_X1 port map( A => net47294, ZN => net56205);
   U39 : INV_X1 port map( A => FUNC(0), ZN => net47294);
   U40 : NAND3_X1 port map( A1 => net56011, A2 => net51772, A3 => net47294, ZN 
                           => net47283);
   U41 : NAND3_X1 port map( A1 => n16, A2 => net47280, A3 => net47281, ZN => 
                           n14);
   U42 : INV_X1 port map( A => net47282, ZN => net47280);
   U43 : AND3_X1 port map( A1 => net54989, A2 => n16, A3 => net47281, ZN => 
                           net54984);
   U44 : NAND2_X1 port map( A1 => n16, A2 => net47281, ZN => net47289);
   U45 : INV_X1 port map( A => FUNC(2), ZN => net47288);
   U46 : INV_X1 port map( A => FUNC(1), ZN => net56055);
   U47 : AOI222_X1 port map( A1 => N63, A2 => net51575, B1 => N95, B2 => 
                           net51581, C1 => Y_LOGIC_16_port, C2 => net51587, ZN 
                           => net47243);
   U48 : BUF_X2 port map( A => n18, Z => net51587);
   U49 : BUF_X2 port map( A => net54984, Z => net51581);
   U50 : BUF_X2 port map( A => n19, Z => net51575);
   U51 : NAND2_X1 port map( A1 => net47283, A2 => net47284, ZN => n18);
   U52 : BUF_X2 port map( A => n18, Z => net51585);
   U53 : BUF_X2 port map( A => net54984, Z => net51583);
   U54 : AND3_X1 port map( A1 => net54989, A2 => net55932, A3 => net51772, ZN 
                           => n19);
   U55 : BUF_X2 port map( A => n19, Z => net51573);
   U56 : BUF_X2 port map( A => n19, Z => net51577);
   U57 : INV_X1 port map( A => n214, ZN => n20);
   U58 : CLKBUF_X1 port map( A => DATA1(13), Z => n21);
   U59 : CLKBUF_X1 port map( A => DATA2(18), Z => n22);
   U60 : INV_X1 port map( A => n219, ZN => n23);
   U61 : CLKBUF_X1 port map( A => DATA2(15), Z => n24);
   U62 : CLKBUF_X1 port map( A => DATA2(26), Z => n25);
   U63 : BUF_X1 port map( A => DATA2(8), Z => n26);
   U64 : INV_X1 port map( A => n244, ZN => n27);
   U65 : INV_X1 port map( A => n248, ZN => n28);
   U66 : INV_X1 port map( A => n247, ZN => n29);
   U67 : INV_X1 port map( A => n245, ZN => n30);
   U68 : INV_X1 port map( A => n225, ZN => n31);
   U69 : INV_X1 port map( A => n204, ZN => n33);
   U70 : CLKBUF_X1 port map( A => DATA1(14), Z => n34);
   U71 : INV_X1 port map( A => n213, ZN => n35);
   U72 : CLKBUF_X1 port map( A => DATA1(0), Z => n36);
   U73 : CLKBUF_X1 port map( A => DATA1(9), Z => n37);
   U74 : INV_X1 port map( A => n211, ZN => n38);
   U75 : INV_X1 port map( A => n253, ZN => n39);
   U76 : CLKBUF_X1 port map( A => DATA1(29), Z => n40);
   U77 : INV_X1 port map( A => n252, ZN => n41);
   U78 : CLKBUF_X1 port map( A => n26, Z => n42);
   U79 : BUF_X2 port map( A => DATA2(1), Z => n43);
   U80 : INV_X1 port map( A => n248, ZN => n44);
   U81 : INV_X1 port map( A => n255, ZN => n45);
   U82 : CLKBUF_X1 port map( A => DATA2(8), Z => n46);
   U83 : INV_X1 port map( A => n256, ZN => n47_port);
   U84 : INV_X1 port map( A => n215, ZN => n48_port);
   U85 : CLKBUF_X1 port map( A => DATA2(22), Z => n49_port);
   U86 : CLKBUF_X1 port map( A => DATA2(3), Z => n50_port);
   U87 : INV_X1 port map( A => n218, ZN => n51_port);
   U88 : BUF_X1 port map( A => n89_port, Z => n113_port);
   U89 : INV_X1 port map( A => n227, ZN => n52_port);
   U90 : CLKBUF_X1 port map( A => DATA1(6), Z => n53_port);
   U91 : CLKBUF_X1 port map( A => DATA2(20), Z => n54_port);
   U92 : INV_X1 port map( A => n223, ZN => n55_port);
   U93 : INV_X1 port map( A => DATA2(0), ZN => n56_port);
   U94 : INV_X2 port map( A => n56_port, ZN => n57_port);
   U95 : INV_X1 port map( A => n208, ZN => n58_port);
   U96 : CLKBUF_X1 port map( A => DATA1(24), Z => n59_port);
   U97 : INV_X1 port map( A => n217, ZN => n60_port);
   U98 : INV_X1 port map( A => n213, ZN => n61_port);
   U99 : CLKBUF_X1 port map( A => DATA2(18), Z => n62_port);
   U100 : CLKBUF_X1 port map( A => DATA2(30), Z => n63_port);
   U101 : INV_X1 port map( A => n205, ZN => n64_port);
   U102 : CLKBUF_X1 port map( A => DATA2(3), Z => n65_port);
   U103 : INV_X1 port map( A => n43, ZN => n66_port);
   U104 : INV_X2 port map( A => n66_port, ZN => n67_port);
   U105 : CLKBUF_X1 port map( A => DATA2(4), Z => n68_port);
   U106 : INV_X1 port map( A => n225, ZN => n69_port);
   U107 : INV_X1 port map( A => n215, ZN => n70_port);
   U108 : CLKBUF_X1 port map( A => DATA2(10), Z => n71_port);
   U109 : CLKBUF_X1 port map( A => DATA2(2), Z => n72_port);
   U110 : INV_X1 port map( A => n212, ZN => n73_port);
   U111 : INV_X1 port map( A => n224, ZN => n74_port);
   U112 : CLKBUF_X1 port map( A => DATA2(11), Z => n75_port);
   U113 : INV_X1 port map( A => n216, ZN => n76_port);
   U114 : NAND2_X1 port map( A1 => N64, A2 => net51573, ZN => n77_port);
   U115 : NAND2_X1 port map( A1 => N96, A2 => net51581, ZN => n78_port);
   U116 : NAND2_X1 port map( A1 => Y_LOGIC_17_port, A2 => net51587, ZN => 
                           n79_port);
   U117 : AND3_X1 port map( A1 => n77_port, A2 => n78_port, A3 => n79_port, ZN 
                           => n170);
   U118 : CLKBUF_X1 port map( A => DATA1(2), Z => n80_port);
   U119 : AND2_X1 port map( A1 => n93_port, A2 => n92_port, ZN => n81_port);
   U120 : AND2_X1 port map( A1 => n91_port, A2 => n81_port, ZN => n152);
   U121 : INV_X1 port map( A => n220, ZN => n82_port);
   U122 : AND2_X1 port map( A1 => n103_port, A2 => n102_port, ZN => n83_port);
   U123 : AND2_X1 port map( A1 => n101_port, A2 => n83_port, ZN => n160);
   U124 : AND2_X1 port map( A1 => n114, A2 => n116, ZN => n84_port);
   U125 : AND2_X1 port map( A1 => n115, A2 => n84_port, ZN => n172);
   U126 : INV_X1 port map( A => n66_port, ZN => n85_port);
   U127 : CLKBUF_X1 port map( A => DATA1(28), Z => n86_port);
   U128 : INV_X1 port map( A => n224, ZN => n87_port);
   U129 : AND2_X1 port map( A1 => n95_port, A2 => n96_port, ZN => n88_port);
   U130 : AND2_X1 port map( A1 => n94_port, A2 => n88_port, ZN => n190);
   U131 : CLKBUF_X1 port map( A => DATA1(8), Z => n89_port);
   U132 : INV_X1 port map( A => n259, ZN => n90_port);
   U133 : NAND2_X1 port map( A1 => N86, A2 => net51579, ZN => n91_port);
   U134 : NAND2_X1 port map( A1 => Y_LOGIC_7_port, A2 => net51585, ZN => 
                           n92_port);
   U135 : NAND2_X1 port map( A1 => N54, A2 => net51577, ZN => n93_port);
   U136 : NAND2_X1 port map( A1 => N74, A2 => net51573, ZN => n94_port);
   U137 : NAND2_X1 port map( A1 => N106, A2 => net51579, ZN => n95_port);
   U138 : NAND2_X1 port map( A1 => Y_LOGIC_27_port, A2 => net51585, ZN => 
                           n96_port);
   U139 : INV_X1 port map( A => n221, ZN => n98_port);
   U140 : INV_X1 port map( A => n257, ZN => n99_port);
   U141 : INV_X1 port map( A => n228, ZN => n100_port);
   U142 : NAND2_X1 port map( A1 => N90, A2 => net51579, ZN => n101_port);
   U143 : NAND2_X1 port map( A1 => Y_LOGIC_11_port, A2 => net51585, ZN => 
                           n102_port);
   U144 : NAND2_X1 port map( A1 => N58, A2 => net51577, ZN => n103_port);
   U145 : NAND2_X1 port map( A1 => N72, A2 => net51573, ZN => n104_port);
   U146 : NAND2_X1 port map( A1 => N104, A2 => net51579, ZN => n105_port);
   U147 : NAND2_X1 port map( A1 => Y_LOGIC_25_port, A2 => net51585, ZN => 
                           n106_port);
   U148 : AND3_X1 port map( A1 => n104_port, A2 => n105_port, A3 => n106_port, 
                           ZN => n186);
   U149 : CLKBUF_X1 port map( A => n57_port, Z => n107_port);
   U150 : NAND2_X1 port map( A1 => N66, A2 => net51573, ZN => n108_port);
   U151 : NAND2_X1 port map( A1 => N98, A2 => net51581, ZN => n109_port);
   U152 : NAND2_X1 port map( A1 => Y_LOGIC_19_port, A2 => net51587, ZN => 
                           n110_port);
   U153 : AND3_X1 port map( A1 => n108_port, A2 => n109_port, A3 => n110_port, 
                           ZN => n174);
   U154 : INV_X1 port map( A => n258, ZN => n111_port);
   U155 : INV_X1 port map( A => n135, ZN => n112_port);
   U156 : NAND2_X1 port map( A1 => N65, A2 => net51573, ZN => n114);
   U157 : NAND2_X1 port map( A1 => N97, A2 => net51581, ZN => n115);
   U158 : NAND2_X1 port map( A1 => Y_LOGIC_18_port, A2 => net51587, ZN => n116)
                           ;
   U159 : NAND2_X1 port map( A1 => N105, A2 => net51579, ZN => n117);
   U160 : NAND2_X1 port map( A1 => Y_LOGIC_26_port, A2 => net51585, ZN => n118)
                           ;
   U161 : NAND2_X1 port map( A1 => N73, A2 => net51577, ZN => n119);
   U162 : AND3_X1 port map( A1 => n117, A2 => n118, A3 => n119, ZN => n188);
   U163 : NAND2_X1 port map( A1 => N101, A2 => net51579, ZN => n120);
   U164 : NAND2_X1 port map( A1 => N69, A2 => net51577, ZN => n121);
   U165 : NAND2_X1 port map( A1 => Y_LOGIC_22_port, A2 => net51587, ZN => n122)
                           ;
   U166 : AND3_X1 port map( A1 => n120, A2 => n121, A3 => n122, ZN => n180);
   U167 : NAND2_X1 port map( A1 => N78, A2 => net51575, ZN => n123);
   U168 : NAND2_X1 port map( A1 => N110, A2 => net51581, ZN => n124);
   U169 : NAND2_X1 port map( A1 => Y_LOGIC_31_port, A2 => net51587, ZN => n125)
                           ;
   U170 : AND3_X1 port map( A1 => n123, A2 => n124, A3 => n125, ZN => n197);
   U171 : NAND2_X1 port map( A1 => N77, A2 => net51573, ZN => n126);
   U172 : NAND2_X1 port map( A1 => N109, A2 => net51579, ZN => n127);
   U173 : NAND2_X1 port map( A1 => Y_LOGIC_30_port, A2 => net51585, ZN => n128)
                           ;
   U174 : AND3_X1 port map( A1 => n126, A2 => n127, A3 => n128, ZN => n195);
   U175 : BUF_X2 port map( A => net23929, Z => net51563);
   U176 : BUF_X2 port map( A => net23929, Z => net51567);
   U177 : BUF_X2 port map( A => net23929, Z => net51565);
   U178 : BUF_X2 port map( A => net23929, Z => net51569);
   U179 : BUF_X2 port map( A => net23929, Z => net51561);
   U180 : BUF_X2 port map( A => S_3_port, Z => n132);
   U181 : BUF_X1 port map( A => S_3_port, Z => n131);
   U182 : BUF_X2 port map( A => S_3_port, Z => n133);
   U183 : CLKBUF_X1 port map( A => DATA1(4), Z => n130);
   U184 : CLKBUF_X1 port map( A => net23929, Z => net51571);
   U185 : INV_X1 port map( A => n107_port, ZN => n134);
   U186 : INV_X1 port map( A => n72_port, ZN => n135);
   U187 : OAI21_X1 port map( B1 => net55932, B2 => net47283, A => net47284, ZN 
                           => S_3_port);
   U188 : INV_X1 port map( A => net47283, ZN => net23929);
   U189 : INV_X1 port map( A => DATA2(31), ZN => n230);
   U190 : INV_X1 port map( A => DATA2(30), ZN => n231);
   U191 : INV_X1 port map( A => DATA2(29), ZN => n232);
   U192 : INV_X1 port map( A => DATA2(28), ZN => n233);
   U193 : INV_X1 port map( A => DATA2(27), ZN => n234);
   U194 : INV_X1 port map( A => DATA2(26), ZN => n235);
   U195 : INV_X1 port map( A => DATA2(25), ZN => n236);
   U196 : INV_X1 port map( A => DATA2(24), ZN => n237);
   U197 : INV_X1 port map( A => DATA2(23), ZN => n238);
   U198 : INV_X1 port map( A => DATA2(22), ZN => n239);
   U199 : INV_X1 port map( A => DATA2(21), ZN => n240);
   U200 : INV_X1 port map( A => DATA2(20), ZN => n241);
   U201 : INV_X1 port map( A => DATA2(19), ZN => n242);
   U202 : INV_X1 port map( A => n22, ZN => n243);
   U203 : INV_X1 port map( A => DATA2(17), ZN => n244);
   U204 : INV_X1 port map( A => DATA2(16), ZN => n245);
   U205 : INV_X1 port map( A => DATA2(15), ZN => n246);
   U206 : INV_X1 port map( A => DATA2(14), ZN => n247);
   U207 : INV_X1 port map( A => DATA2(13), ZN => n248);
   U208 : INV_X1 port map( A => DATA2(12), ZN => n249);
   U209 : INV_X1 port map( A => DATA2(11), ZN => n250);
   U210 : INV_X1 port map( A => DATA2(10), ZN => n251);
   U211 : INV_X1 port map( A => DATA2(9), ZN => n252);
   U212 : INV_X1 port map( A => n42, ZN => n253);
   U213 : INV_X1 port map( A => DATA2(7), ZN => n254);
   U214 : INV_X1 port map( A => DATA2(6), ZN => n255);
   U215 : INV_X1 port map( A => DATA2(5), ZN => n256);
   U216 : INV_X1 port map( A => n68_port, ZN => n257);
   U217 : INV_X1 port map( A => n65_port, ZN => n258);
   U218 : INV_X1 port map( A => DATA1(31), ZN => n199);
   U219 : INV_X1 port map( A => DATA1(30), ZN => n200);
   U220 : INV_X1 port map( A => DATA1(29), ZN => n201);
   U221 : INV_X1 port map( A => n86_port, ZN => n202);
   U222 : INV_X1 port map( A => DATA1(27), ZN => n203);
   U223 : INV_X1 port map( A => DATA1(26), ZN => n204);
   U224 : INV_X1 port map( A => DATA1(25), ZN => n205);
   U225 : INV_X1 port map( A => DATA1(24), ZN => n206);
   U226 : INV_X1 port map( A => DATA1(23), ZN => n207);
   U227 : INV_X1 port map( A => DATA1(22), ZN => n208);
   U228 : INV_X1 port map( A => DATA1(21), ZN => n209);
   U229 : INV_X1 port map( A => DATA1(20), ZN => n210);
   U230 : INV_X1 port map( A => DATA1(19), ZN => n211);
   U231 : INV_X1 port map( A => DATA1(18), ZN => n212);
   U232 : INV_X1 port map( A => DATA1(17), ZN => n213);
   U233 : INV_X1 port map( A => DATA1(16), ZN => n214);
   U234 : INV_X1 port map( A => DATA1(15), ZN => n215);
   U235 : INV_X1 port map( A => DATA1(14), ZN => n216);
   U236 : INV_X1 port map( A => n21, ZN => n217);
   U237 : INV_X1 port map( A => DATA1(12), ZN => n218);
   U238 : INV_X1 port map( A => DATA1(11), ZN => n219);
   U239 : INV_X1 port map( A => DATA1(10), ZN => n220);
   U240 : INV_X1 port map( A => n37, ZN => n221);
   U241 : INV_X1 port map( A => n113_port, ZN => n222);
   U242 : INV_X1 port map( A => DATA1(7), ZN => n223);
   U243 : INV_X1 port map( A => DATA1(6), ZN => n224);
   U244 : INV_X1 port map( A => DATA1(5), ZN => n225);
   U245 : INV_X1 port map( A => DATA1(4), ZN => n226);
   U246 : INV_X1 port map( A => DATA1(3), ZN => n227);
   U247 : INV_X1 port map( A => n80_port, ZN => n228);
   U248 : INV_X1 port map( A => n129, ZN => n229);
   U249 : INV_X1 port map( A => n36, ZN => n259);
   U250 : NAND2_X1 port map( A1 => N113, A2 => net51772, ZN => net47291);
   U251 : OAI221_X1 port map( B1 => N112, B2 => net47281, C1 => N111, C2 => 
                           net47289, A => net47290, ZN => n139);
   U252 : NAND2_X1 port map( A1 => N47, A2 => net51577, ZN => n138);
   U253 : AOI22_X1 port map( A1 => N79, A2 => net51579, B1 => Y_LOGIC_0_port, 
                           B2 => net51585, ZN => n137);
   U254 : NAND2_X1 port map( A1 => OUT_SHIFTER_0_port, A2 => net51591, ZN => 
                           n136);
   U255 : NAND4_X1 port map( A1 => n136, A2 => n138, A3 => n137, A4 => n139, ZN
                           => OUTALU(0));
   U256 : NAND2_X1 port map( A1 => OUT_SHIFTER_1_port, A2 => net51591, ZN => 
                           n141);
   U257 : AOI222_X1 port map( A1 => N48, A2 => net51577, B1 => N80, B2 => 
                           net51579, C1 => Y_LOGIC_1_port, C2 => net51585, ZN 
                           => n140);
   U258 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => OUTALU(1));
   U259 : NAND2_X1 port map( A1 => OUT_SHIFTER_2_port, A2 => net51591, ZN => 
                           n143);
   U260 : AOI222_X1 port map( A1 => N49, A2 => net51577, B1 => N81, B2 => 
                           net51583, C1 => Y_LOGIC_2_port, C2 => net51589, ZN 
                           => n142);
   U261 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => OUTALU(2));
   U262 : NAND2_X1 port map( A1 => OUT_SHIFTER_3_port, A2 => net51591, ZN => 
                           n145);
   U263 : AOI222_X1 port map( A1 => N50, A2 => net51575, B1 => N82, B2 => 
                           net51583, C1 => Y_LOGIC_3_port, C2 => net51589, ZN 
                           => n144);
   U264 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => OUTALU(3));
   U265 : NAND2_X1 port map( A1 => OUT_SHIFTER_4_port, A2 => net51591, ZN => 
                           n147);
   U266 : AOI222_X1 port map( A1 => N51, A2 => net51577, B1 => N83, B2 => 
                           net51583, C1 => Y_LOGIC_4_port, C2 => net51589, ZN 
                           => n146);
   U267 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => OUTALU(4));
   U268 : NAND2_X1 port map( A1 => OUT_SHIFTER_5_port, A2 => net51591, ZN => 
                           n149);
   U269 : AOI222_X1 port map( A1 => N52, A2 => net51575, B1 => N84, B2 => 
                           net51583, C1 => Y_LOGIC_5_port, C2 => net51589, ZN 
                           => n148);
   U270 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => OUTALU(5));
   U271 : NAND2_X1 port map( A1 => OUT_SHIFTER_6_port, A2 => net51591, ZN => 
                           n151);
   U272 : AOI222_X1 port map( A1 => N53, A2 => net51575, B1 => N85, B2 => 
                           net51583, C1 => Y_LOGIC_6_port, C2 => net51589, ZN 
                           => n150);
   U273 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => OUTALU(6));
   U274 : NAND2_X1 port map( A1 => OUT_SHIFTER_7_port, A2 => net51591, ZN => 
                           n153);
   U275 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => OUTALU(7));
   U276 : NAND2_X1 port map( A1 => OUT_SHIFTER_8_port, A2 => net51591, ZN => 
                           n155);
   U277 : AOI222_X1 port map( A1 => N55, A2 => net51575, B1 => N87, B2 => 
                           net51583, C1 => Y_LOGIC_8_port, C2 => net51589, ZN 
                           => n154);
   U278 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => OUTALU(8));
   U279 : NAND2_X1 port map( A1 => OUT_SHIFTER_9_port, A2 => net51591, ZN => 
                           n157);
   U280 : AOI222_X1 port map( A1 => N56, A2 => net51575, B1 => N88, B2 => 
                           net51583, C1 => Y_LOGIC_9_port, C2 => net51589, ZN 
                           => n156);
   U281 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => OUTALU(9));
   U282 : NAND2_X1 port map( A1 => OUT_SHIFTER_10_port, A2 => net51591, ZN => 
                           n159);
   U283 : AOI222_X1 port map( A1 => N57, A2 => net51575, B1 => N89, B2 => 
                           net51583, C1 => Y_LOGIC_10_port, C2 => net51589, ZN 
                           => n158);
   U284 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => OUTALU(10));
   U285 : NAND2_X1 port map( A1 => OUT_SHIFTER_11_port, A2 => net51591, ZN => 
                           n161);
   U286 : NAND2_X1 port map( A1 => n161, A2 => n160, ZN => OUTALU(11));
   U287 : NAND2_X1 port map( A1 => OUT_SHIFTER_12_port, A2 => net51593, ZN => 
                           n163);
   U288 : AOI222_X1 port map( A1 => N59, A2 => net51575, B1 => N91, B2 => 
                           net51581, C1 => Y_LOGIC_12_port, C2 => net51587, ZN 
                           => n162);
   U289 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => OUTALU(12));
   U290 : NAND2_X1 port map( A1 => OUT_SHIFTER_13_port, A2 => net51593, ZN => 
                           n165);
   U291 : AOI222_X1 port map( A1 => N60, A2 => net51575, B1 => N92, B2 => 
                           net51581, C1 => Y_LOGIC_13_port, C2 => net51587, ZN 
                           => n164);
   U292 : NAND2_X1 port map( A1 => n165, A2 => n164, ZN => OUTALU(13));
   U293 : NAND2_X1 port map( A1 => OUT_SHIFTER_14_port, A2 => net51593, ZN => 
                           n167);
   U294 : AOI222_X1 port map( A1 => N61, A2 => net51575, B1 => N93, B2 => 
                           net51581, C1 => Y_LOGIC_14_port, C2 => net51587, ZN 
                           => n166);
   U295 : NAND2_X1 port map( A1 => n167, A2 => n166, ZN => OUTALU(14));
   U296 : NAND2_X1 port map( A1 => OUT_SHIFTER_15_port, A2 => net51593, ZN => 
                           n169);
   U297 : AOI222_X1 port map( A1 => N62, A2 => net51575, B1 => N94, B2 => 
                           net51581, C1 => Y_LOGIC_15_port, C2 => net51587, ZN 
                           => n168);
   U298 : NAND2_X1 port map( A1 => n169, A2 => n168, ZN => OUTALU(15));
   U299 : NAND2_X1 port map( A1 => OUT_SHIFTER_17_port, A2 => net51593, ZN => 
                           n171);
   U300 : NAND2_X1 port map( A1 => n171, A2 => n170, ZN => OUTALU(17));
   U301 : NAND2_X1 port map( A1 => OUT_SHIFTER_18_port, A2 => net51593, ZN => 
                           n173);
   U302 : NAND2_X1 port map( A1 => n173, A2 => n172, ZN => OUTALU(18));
   U303 : NAND2_X1 port map( A1 => OUT_SHIFTER_19_port, A2 => net51593, ZN => 
                           n175);
   U304 : NAND2_X1 port map( A1 => n175, A2 => n174, ZN => OUTALU(19));
   U305 : NAND2_X1 port map( A1 => OUT_SHIFTER_20_port, A2 => net51593, ZN => 
                           n177);
   U306 : AOI222_X1 port map( A1 => N67, A2 => net51573, B1 => N99, B2 => 
                           net51581, C1 => Y_LOGIC_20_port, C2 => net51587, ZN 
                           => n176);
   U307 : NAND2_X1 port map( A1 => n177, A2 => n176, ZN => OUTALU(20));
   U308 : NAND2_X1 port map( A1 => OUT_SHIFTER_21_port, A2 => net51593, ZN => 
                           n179);
   U309 : AOI222_X1 port map( A1 => N68, A2 => net51573, B1 => N100, B2 => 
                           net51581, C1 => Y_LOGIC_21_port, C2 => net51587, ZN 
                           => n178);
   U310 : NAND2_X1 port map( A1 => n179, A2 => n178, ZN => OUTALU(21));
   U311 : NAND2_X1 port map( A1 => OUT_SHIFTER_22_port, A2 => net51593, ZN => 
                           n181);
   U312 : NAND2_X1 port map( A1 => n181, A2 => n180, ZN => OUTALU(22));
   U313 : NAND2_X1 port map( A1 => OUT_SHIFTER_23_port, A2 => net51593, ZN => 
                           n183);
   U314 : AOI222_X1 port map( A1 => N70, A2 => net51573, B1 => N102, B2 => 
                           net51581, C1 => Y_LOGIC_23_port, C2 => net51585, ZN 
                           => n182);
   U315 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => OUTALU(23));
   U316 : NAND2_X1 port map( A1 => OUT_SHIFTER_24_port, A2 => net51595, ZN => 
                           n185);
   U317 : AOI222_X1 port map( A1 => N71, A2 => net51573, B1 => N103, B2 => 
                           net51579, C1 => Y_LOGIC_24_port, C2 => net51585, ZN 
                           => n184);
   U318 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => OUTALU(24));
   U319 : NAND2_X1 port map( A1 => OUT_SHIFTER_25_port, A2 => net51595, ZN => 
                           n187);
   U320 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => OUTALU(25));
   U321 : NAND2_X1 port map( A1 => OUT_SHIFTER_26_port, A2 => net51595, ZN => 
                           n189);
   U322 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => OUTALU(26));
   U323 : NAND2_X1 port map( A1 => OUT_SHIFTER_27_port, A2 => net51595, ZN => 
                           n191);
   U324 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => OUTALU(27));
   U325 : NAND2_X1 port map( A1 => OUT_SHIFTER_28_port, A2 => net51595, ZN => 
                           n192);
   U326 : NAND2_X1 port map( A1 => n192, A2 => n3, ZN => OUTALU(28));
   U327 : NAND2_X1 port map( A1 => OUT_SHIFTER_29_port, A2 => net51595, ZN => 
                           n194);
   U328 : AOI222_X1 port map( A1 => N76, A2 => net51573, B1 => N108, B2 => 
                           net51579, C1 => Y_LOGIC_29_port, C2 => net51585, ZN 
                           => n193);
   U329 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => OUTALU(29));
   U330 : NAND2_X1 port map( A1 => net51595, A2 => OUT_SHIFTER_30_port, ZN => 
                           n196);
   U331 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => OUTALU(30));
   U332 : NAND2_X1 port map( A1 => OUT_SHIFTER_31_port, A2 => net51595, ZN => 
                           n198);
   U333 : NAND2_X1 port map( A1 => n197, A2 => n198, ZN => OUTALU(31));
   NAND31I_1 : NAND3_0 port map( A => n259, B => n134, C => X_Logic0_port, Y =>
                           L0_0_port);
   NAND31I_2 : NAND3_127 port map( A => n229, B => n66_port, C => X_Logic0_port
                           , Y => L0_1_port);
   NAND31I_3 : NAND3_126 port map( A => n228, B => n135, C => X_Logic0_port, Y 
                           => L0_2_port);
   NAND31I_4 : NAND3_125 port map( A => n227, B => n258, C => X_Logic0_port, Y 
                           => L0_3_port);
   NAND31I_5 : NAND3_124 port map( A => n226, B => n257, C => X_Logic0_port, Y 
                           => L0_4_port);
   NAND31I_6 : NAND3_123 port map( A => n225, B => n256, C => X_Logic0_port, Y 
                           => L0_5_port);
   NAND31I_7 : NAND3_122 port map( A => n224, B => n255, C => X_Logic0_port, Y 
                           => L0_6_port);
   NAND31I_8 : NAND3_121 port map( A => n223, B => n254, C => X_Logic0_port, Y 
                           => L0_7_port);
   NAND31I_9 : NAND3_120 port map( A => n222, B => n253, C => X_Logic0_port, Y 
                           => L0_8_port);
   NAND31I_10 : NAND3_119 port map( A => n221, B => n252, C => X_Logic0_port, Y
                           => L0_9_port);
   NAND31I_11 : NAND3_118 port map( A => n220, B => n251, C => X_Logic0_port, Y
                           => L0_10_port);
   NAND31I_12 : NAND3_117 port map( A => n219, B => n250, C => X_Logic0_port, Y
                           => L0_11_port);
   NAND31I_13 : NAND3_116 port map( A => n218, B => n249, C => X_Logic0_port, Y
                           => L0_12_port);
   NAND31I_14 : NAND3_115 port map( A => n217, B => n248, C => X_Logic0_port, Y
                           => L0_13_port);
   NAND31I_15 : NAND3_114 port map( A => n216, B => n247, C => X_Logic0_port, Y
                           => L0_14_port);
   NAND31I_16 : NAND3_113 port map( A => n215, B => n246, C => X_Logic0_port, Y
                           => L0_15_port);
   NAND31I_17 : NAND3_112 port map( A => n214, B => n245, C => X_Logic0_port, Y
                           => L0_16_port);
   NAND31I_18 : NAND3_111 port map( A => n213, B => n244, C => X_Logic0_port, Y
                           => L0_17_port);
   NAND31I_19 : NAND3_110 port map( A => n212, B => n243, C => X_Logic0_port, Y
                           => L0_18_port);
   NAND31I_20 : NAND3_109 port map( A => n211, B => n242, C => X_Logic0_port, Y
                           => L0_19_port);
   NAND31I_21 : NAND3_108 port map( A => n210, B => n241, C => X_Logic0_port, Y
                           => L0_20_port);
   NAND31I_22 : NAND3_107 port map( A => n209, B => n240, C => X_Logic0_port, Y
                           => L0_21_port);
   NAND31I_23 : NAND3_106 port map( A => n208, B => n239, C => X_Logic0_port, Y
                           => L0_22_port);
   NAND31I_24 : NAND3_105 port map( A => n207, B => n238, C => X_Logic0_port, Y
                           => L0_23_port);
   NAND31I_25 : NAND3_104 port map( A => n206, B => n237, C => X_Logic0_port, Y
                           => L0_24_port);
   NAND31I_26 : NAND3_103 port map( A => n205, B => n236, C => X_Logic0_port, Y
                           => L0_25_port);
   NAND31I_27 : NAND3_102 port map( A => n204, B => n235, C => X_Logic0_port, Y
                           => L0_26_port);
   NAND31I_28 : NAND3_101 port map( A => n203, B => n234, C => X_Logic0_port, Y
                           => L0_27_port);
   NAND31I_29 : NAND3_100 port map( A => n202, B => n233, C => X_Logic0_port, Y
                           => L0_28_port);
   NAND31I_30 : NAND3_99 port map( A => n201, B => n232, C => X_Logic0_port, Y 
                           => L0_29_port);
   NAND31I_31 : NAND3_98 port map( A => n200, B => n231, C => X_Logic0_port, Y 
                           => L0_30_port);
   NAND31I_32 : NAND3_97 port map( A => n199, B => n230, C => X_Logic0_port, Y 
                           => L0_31_port);
   NAND31I_1_0 : NAND3_96 port map( A => n259, B => n107_port, C => net51561, Y
                           => L1_0_port);
   NAND31I_2_0 : NAND3_95 port map( A => n229, B => n85_port, C => net51561, Y 
                           => L1_1_port);
   NAND31I_3_0 : NAND3_94 port map( A => n228, B => n112_port, C => net51561, Y
                           => L1_2_port);
   NAND31I_4_0 : NAND3_93 port map( A => n227, B => n111_port, C => net51561, Y
                           => L1_3_port);
   NAND31I_5_0 : NAND3_92 port map( A => n226, B => n68_port, C => net51561, Y 
                           => L1_4_port);
   NAND31I_6_0 : NAND3_91 port map( A => n225, B => n47_port, C => net51561, Y 
                           => L1_5_port);
   NAND31I_7_0 : NAND3_90 port map( A => n224, B => n45, C => net51561, Y => 
                           L1_6_port);
   NAND31I_8_0 : NAND3_89 port map( A => n223, B => DATA2(7), C => net51561, Y 
                           => L1_7_port);
   NAND31I_9_0 : NAND3_88 port map( A => n222, B => n46, C => net51561, Y => 
                           L1_8_port);
   NAND31I_10_0 : NAND3_87 port map( A => n221, B => n41, C => net51561, Y => 
                           L1_9_port);
   NAND31I_11_0 : NAND3_86 port map( A => n220, B => n71_port, C => net51561, Y
                           => L1_10_port);
   NAND31I_12_0 : NAND3_85 port map( A => n219, B => n75_port, C => net51561, Y
                           => L1_11_port);
   NAND31I_13_0 : NAND3_84 port map( A => n218, B => DATA2(12), C => net51563, 
                           Y => L1_12_port);
   NAND31I_14_0 : NAND3_83 port map( A => n217, B => n44, C => net51563, Y => 
                           L1_13_port);
   NAND31I_15_0 : NAND3_82 port map( A => n216, B => n29, C => net51563, Y => 
                           L1_14_port);
   NAND31I_16_0 : NAND3_81 port map( A => n215, B => n24, C => net51563, Y => 
                           L1_15_port);
   NAND31I_17_0 : NAND3_80 port map( A => n214, B => n30, C => net51563, Y => 
                           L1_16_port);
   NAND31I_18_0 : NAND3_79 port map( A => n213, B => n27, C => net51563, Y => 
                           L1_17_port);
   NAND31I_19_0 : NAND3_78 port map( A => n212, B => n62_port, C => net51563, Y
                           => L1_18_port);
   NAND31I_20_0 : NAND3_77 port map( A => n211, B => DATA2(19), C => net51563, 
                           Y => L1_19_port);
   NAND31I_21_0 : NAND3_76 port map( A => n210, B => n54_port, C => net51563, Y
                           => L1_20_port);
   NAND31I_22_0 : NAND3_75 port map( A => n209, B => DATA2(21), C => net51563, 
                           Y => L1_21_port);
   NAND31I_23_0 : NAND3_74 port map( A => n208, B => n49_port, C => net51563, Y
                           => L1_22_port);
   NAND31I_24_0 : NAND3_73 port map( A => n207, B => DATA2(23), C => net51563, 
                           Y => L1_23_port);
   NAND31I_25_0 : NAND3_72 port map( A => n206, B => DATA2(24), C => net51565, 
                           Y => L1_24_port);
   NAND31I_26_0 : NAND3_71 port map( A => n205, B => DATA2(25), C => net51565, 
                           Y => L1_25_port);
   NAND31I_27_0 : NAND3_70 port map( A => n204, B => n25, C => net51565, Y => 
                           L1_26_port);
   NAND31I_28_0 : NAND3_69 port map( A => n203, B => DATA2(27), C => net51565, 
                           Y => L1_27_port);
   NAND31I_29_0 : NAND3_68 port map( A => n202, B => DATA2(28), C => net51565, 
                           Y => L1_28_port);
   NAND31I_30_0 : NAND3_67 port map( A => n201, B => DATA2(29), C => net51565, 
                           Y => L1_29_port);
   NAND31I_31_0 : NAND3_66 port map( A => n200, B => n63_port, C => net51565, Y
                           => L1_30_port);
   NAND31I_32_0 : NAND3_65 port map( A => n199, B => DATA2(31), C => net51565, 
                           Y => L1_31_port);
   NAND31I_1_1 : NAND3_64 port map( A => n90_port, B => n134, C => net51565, Y 
                           => L2_0_port);
   NAND31I_2_1 : NAND3_63 port map( A => n129, B => n66_port, C => net51565, Y 
                           => L2_1_port);
   NAND31I_3_1 : NAND3_62 port map( A => n100_port, B => n135, C => net51565, Y
                           => L2_2_port);
   NAND31I_4_1 : NAND3_61 port map( A => n52_port, B => n258, C => net51565, Y 
                           => L2_3_port);
   NAND31I_5_1 : NAND3_60 port map( A => n130, B => n257, C => net51567, Y => 
                           L2_4_port);
   NAND31I_6_1 : NAND3_59 port map( A => n69_port, B => n256, C => net51567, Y 
                           => L2_5_port);
   NAND31I_7_1 : NAND3_58 port map( A => n87_port, B => n255, C => net51567, Y 
                           => L2_6_port);
   NAND31I_8_1 : NAND3_57 port map( A => n55_port, B => n254, C => net51567, Y 
                           => L2_7_port);
   NAND31I_9_1 : NAND3_56 port map( A => n113_port, B => n253, C => net51567, Y
                           => L2_8_port);
   NAND31I_10_1 : NAND3_55 port map( A => n98_port, B => n252, C => net51567, Y
                           => L2_9_port);
   NAND31I_11_1 : NAND3_54 port map( A => n82_port, B => n251, C => net51567, Y
                           => L2_10_port);
   NAND31I_12_1 : NAND3_53 port map( A => n23, B => n250, C => net51567, Y => 
                           L2_11_port);
   NAND31I_13_1 : NAND3_52 port map( A => n51_port, B => n249, C => net51567, Y
                           => L2_12_port);
   NAND31I_14_1 : NAND3_51 port map( A => n32, B => n248, C => net51567, Y => 
                           L2_13_port);
   NAND31I_15_1 : NAND3_50 port map( A => n76_port, B => n247, C => net51567, Y
                           => L2_14_port);
   NAND31I_16_1 : NAND3_49 port map( A => n70_port, B => n246, C => net51567, Y
                           => L2_15_port);
   NAND31I_17_1 : NAND3_48 port map( A => n20, B => n245, C => net51569, Y => 
                           L2_16_port);
   NAND31I_18_1 : NAND3_47 port map( A => n61_port, B => n244, C => net51569, Y
                           => L2_17_port);
   NAND31I_19_1 : NAND3_46 port map( A => n73_port, B => n243, C => net51569, Y
                           => L2_18_port);
   NAND31I_20_1 : NAND3_45 port map( A => n38, B => n242, C => net51569, Y => 
                           L2_19_port);
   NAND31I_21_1 : NAND3_44 port map( A => DATA1(20), B => n241, C => net51569, 
                           Y => L2_20_port);
   NAND31I_22_1 : NAND3_43 port map( A => DATA1(21), B => n240, C => net51569, 
                           Y => L2_21_port);
   NAND31I_23_1 : NAND3_42 port map( A => n58_port, B => n239, C => net51569, Y
                           => L2_22_port);
   NAND31I_24_1 : NAND3_41 port map( A => DATA1(23), B => n238, C => net51569, 
                           Y => L2_23_port);
   NAND31I_25_1 : NAND3_40 port map( A => n59_port, B => n237, C => net51569, Y
                           => L2_24_port);
   NAND31I_26_1 : NAND3_39 port map( A => n64_port, B => n236, C => net51569, Y
                           => L2_25_port);
   NAND31I_27_1 : NAND3_38 port map( A => n33, B => n235, C => net51569, Y => 
                           L2_26_port);
   NAND31I_28_1 : NAND3_37 port map( A => DATA1(27), B => n234, C => net51569, 
                           Y => L2_27_port);
   NAND31I_29_1 : NAND3_36 port map( A => n86_port, B => n233, C => net51571, Y
                           => L2_28_port);
   NAND31I_30_1 : NAND3_35 port map( A => n40, B => n232, C => net51571, Y => 
                           L2_29_port);
   NAND31I_31_1 : NAND3_34 port map( A => DATA1(30), B => n231, C => net51571, 
                           Y => L2_30_port);
   NAND31I_32_1 : NAND3_33 port map( A => DATA1(31), B => n230, C => net51571, 
                           Y => L2_31_port);
   NAND31I_1_2 : NAND3_32 port map( A => n90_port, B => n107_port, C => n131, Y
                           => L3_0_port);
   NAND31I_2_2 : NAND3_31 port map( A => n129, B => n85_port, C => n131, Y => 
                           L3_1_port);
   NAND31I_3_2 : NAND3_30 port map( A => n100_port, B => n112_port, C => n131, 
                           Y => L3_2_port);
   NAND31I_4_2 : NAND3_29 port map( A => n52_port, B => n111_port, C => n131, Y
                           => L3_3_port);
   NAND31I_5_2 : NAND3_28 port map( A => n1, B => n99_port, C => n131, Y => 
                           L3_4_port);
   NAND31I_6_2 : NAND3_27 port map( A => n69_port, B => n47_port, C => n131, Y 
                           => L3_5_port);
   NAND31I_7_2 : NAND3_26 port map( A => n53_port, B => n45, C => n131, Y => 
                           L3_6_port);
   NAND31I_8_2 : NAND3_25 port map( A => n55_port, B => DATA2(7), C => n131, Y 
                           => L3_7_port);
   NAND31I_9_2 : NAND3_24 port map( A => n113_port, B => n46, C => n131, Y => 
                           L3_8_port);
   NAND31I_10_2 : NAND3_23 port map( A => n98_port, B => n41, C => n131, Y => 
                           L3_9_port);
   NAND31I_11_2 : NAND3_22 port map( A => n82_port, B => n71_port, C => n131, Y
                           => L3_10_port);
   NAND31I_12_2 : NAND3_21 port map( A => n23, B => n75_port, C => n131, Y => 
                           L3_11_port);
   NAND31I_13_2 : NAND3_20 port map( A => n51_port, B => DATA2(12), C => n132, 
                           Y => L3_12_port);
   NAND31I_14_2 : NAND3_19 port map( A => n32, B => n44, C => n132, Y => 
                           L3_13_port);
   NAND31I_15_2 : NAND3_18 port map( A => n76_port, B => n29, C => n132, Y => 
                           L3_14_port);
   NAND31I_16_2 : NAND3_17 port map( A => n70_port, B => DATA2(15), C => n132, 
                           Y => L3_15_port);
   NAND31I_17_2 : NAND3_16 port map( A => n20, B => n30, C => n132, Y => 
                           L3_16_port);
   NAND31I_18_2 : NAND3_15 port map( A => n61_port, B => n27, C => n132, Y => 
                           L3_17_port);
   NAND31I_19_2 : NAND3_14 port map( A => n73_port, B => n62_port, C => n132, Y
                           => L3_18_port);
   NAND31I_20_2 : NAND3_13 port map( A => n38, B => DATA2(19), C => n132, Y => 
                           L3_19_port);
   NAND31I_21_2 : NAND3_12 port map( A => DATA1(20), B => n54_port, C => n132, 
                           Y => L3_20_port);
   NAND31I_22_2 : NAND3_11 port map( A => DATA1(21), B => DATA2(21), C => n132,
                           Y => L3_21_port);
   NAND31I_23_2 : NAND3_10 port map( A => n58_port, B => n49_port, C => n132, Y
                           => L3_22_port);
   NAND31I_24_2 : NAND3_9 port map( A => DATA1(23), B => DATA2(23), C => n132, 
                           Y => L3_23_port);
   NAND31I_25_2 : NAND3_8 port map( A => n59_port, B => DATA2(24), C => n133, Y
                           => L3_24_port);
   NAND31I_26_2 : NAND3_7 port map( A => DATA1(25), B => DATA2(25), C => n133, 
                           Y => L3_25_port);
   NAND31I_27_2 : NAND3_6 port map( A => DATA1(26), B => n25, C => n133, Y => 
                           L3_26_port);
   NAND31I_28_2 : NAND3_5 port map( A => DATA1(27), B => DATA2(27), C => n133, 
                           Y => L3_27_port);
   NAND31I_29_2 : NAND3_4 port map( A => n86_port, B => DATA2(28), C => n133, Y
                           => L3_28_port);
   NAND31I_30_2 : NAND3_3 port map( A => n40, B => DATA2(29), C => n133, Y => 
                           L3_29_port);
   NAND31I_31_2 : NAND3_2 port map( A => DATA1(30), B => n63_port, C => n133, Y
                           => L3_30_port);
   NAND31I_32_2 : NAND3_1 port map( A => DATA1(31), B => DATA2(31), C => n133, 
                           Y => L3_31_port);
   NAND41I_1 : NAND4_0 port map( A => L0_0_port, B => L1_0_port, C => L2_0_port
                           , D => L3_0_port, Y => Y_LOGIC_0_port);
   NAND41I_2 : NAND4_31 port map( A => L0_1_port, B => L1_1_port, C => 
                           L2_1_port, D => L3_1_port, Y => Y_LOGIC_1_port);
   NAND41I_3 : NAND4_30 port map( A => L0_2_port, B => L1_2_port, C => 
                           L2_2_port, D => L3_2_port, Y => Y_LOGIC_2_port);
   NAND41I_4 : NAND4_29 port map( A => L0_3_port, B => L1_3_port, C => 
                           L2_3_port, D => L3_3_port, Y => Y_LOGIC_3_port);
   NAND41I_5 : NAND4_28 port map( A => L0_4_port, B => L1_4_port, C => 
                           L2_4_port, D => L3_4_port, Y => Y_LOGIC_4_port);
   NAND41I_6 : NAND4_27 port map( A => L0_5_port, B => L1_5_port, C => 
                           L2_5_port, D => L3_5_port, Y => Y_LOGIC_5_port);
   NAND41I_7 : NAND4_26 port map( A => L0_6_port, B => L1_6_port, C => 
                           L2_6_port, D => L3_6_port, Y => Y_LOGIC_6_port);
   NAND41I_8 : NAND4_25 port map( A => L0_7_port, B => L1_7_port, C => 
                           L2_7_port, D => L3_7_port, Y => Y_LOGIC_7_port);
   NAND41I_9 : NAND4_24 port map( A => L0_8_port, B => L1_8_port, C => 
                           L2_8_port, D => L3_8_port, Y => Y_LOGIC_8_port);
   NAND41I_10 : NAND4_23 port map( A => L0_9_port, B => L1_9_port, C => 
                           L2_9_port, D => L3_9_port, Y => Y_LOGIC_9_port);
   NAND41I_11 : NAND4_22 port map( A => L0_10_port, B => L1_10_port, C => 
                           L2_10_port, D => L3_10_port, Y => Y_LOGIC_10_port);
   NAND41I_12 : NAND4_21 port map( A => L0_11_port, B => L1_11_port, C => 
                           L2_11_port, D => L3_11_port, Y => Y_LOGIC_11_port);
   NAND41I_13 : NAND4_20 port map( A => L0_12_port, B => L1_12_port, C => 
                           L2_12_port, D => L3_12_port, Y => Y_LOGIC_12_port);
   NAND41I_14 : NAND4_19 port map( A => L0_13_port, B => L1_13_port, C => 
                           L2_13_port, D => L3_13_port, Y => Y_LOGIC_13_port);
   NAND41I_15 : NAND4_18 port map( A => L0_14_port, B => L1_14_port, C => 
                           L2_14_port, D => L3_14_port, Y => Y_LOGIC_14_port);
   NAND41I_16 : NAND4_17 port map( A => L0_15_port, B => L1_15_port, C => 
                           L2_15_port, D => L3_15_port, Y => Y_LOGIC_15_port);
   NAND41I_17 : NAND4_16 port map( A => L0_16_port, B => L1_16_port, C => 
                           L2_16_port, D => L3_16_port, Y => Y_LOGIC_16_port);
   NAND41I_18 : NAND4_15 port map( A => L0_17_port, B => L1_17_port, C => 
                           L2_17_port, D => L3_17_port, Y => Y_LOGIC_17_port);
   NAND41I_19 : NAND4_14 port map( A => L0_18_port, B => L1_18_port, C => 
                           L2_18_port, D => L3_18_port, Y => Y_LOGIC_18_port);
   NAND41I_20 : NAND4_13 port map( A => L0_19_port, B => L1_19_port, C => 
                           L2_19_port, D => L3_19_port, Y => Y_LOGIC_19_port);
   NAND41I_21 : NAND4_12 port map( A => L0_20_port, B => L1_20_port, C => 
                           L2_20_port, D => L3_20_port, Y => Y_LOGIC_20_port);
   NAND41I_22 : NAND4_11 port map( A => L0_21_port, B => L1_21_port, C => 
                           L2_21_port, D => L3_21_port, Y => Y_LOGIC_21_port);
   NAND41I_23 : NAND4_10 port map( A => L0_22_port, B => L1_22_port, C => 
                           L2_22_port, D => L3_22_port, Y => Y_LOGIC_22_port);
   NAND41I_24 : NAND4_9 port map( A => L0_23_port, B => L1_23_port, C => 
                           L2_23_port, D => L3_23_port, Y => Y_LOGIC_23_port);
   NAND41I_25 : NAND4_8 port map( A => L0_24_port, B => L1_24_port, C => 
                           L2_24_port, D => L3_24_port, Y => Y_LOGIC_24_port);
   NAND41I_26 : NAND4_7 port map( A => L0_25_port, B => L1_25_port, C => 
                           L2_25_port, D => L3_25_port, Y => Y_LOGIC_25_port);
   NAND41I_27 : NAND4_6 port map( A => L0_26_port, B => L1_26_port, C => 
                           L2_26_port, D => L3_26_port, Y => Y_LOGIC_26_port);
   NAND41I_28 : NAND4_5 port map( A => L0_27_port, B => L1_27_port, C => 
                           L2_27_port, D => L3_27_port, Y => Y_LOGIC_27_port);
   NAND41I_29 : NAND4_4 port map( A => L0_28_port, B => L1_28_port, C => 
                           L2_28_port, D => L3_28_port, Y => Y_LOGIC_28_port);
   NAND41I_30 : NAND4_3 port map( A => L0_29_port, B => L1_29_port, C => 
                           L2_29_port, D => L3_29_port, Y => Y_LOGIC_29_port);
   NAND41I_31 : NAND4_2 port map( A => L0_30_port, B => L1_30_port, C => 
                           L2_30_port, D => L3_30_port, Y => Y_LOGIC_30_port);
   NAND41I_32 : NAND4_1 port map( A => L0_31_port, B => L1_31_port, C => 
                           L2_31_port, D => L3_31_port, Y => Y_LOGIC_31_port);
   SHIFTER : BARREL_SHIFTER_N32 port map( CONF => net55526, DATA1(31) => 
                           DATA1(31), DATA1(30) => DATA1(30), DATA1(29) => 
                           DATA1(29), DATA1(28) => DATA1(28), DATA1(27) => 
                           DATA1(27), DATA1(26) => n33, DATA1(25) => n64_port, 
                           DATA1(24) => DATA1(24), DATA1(23) => DATA1(23), 
                           DATA1(22) => DATA1(22), DATA1(21) => DATA1(21), 
                           DATA1(20) => DATA1(20), DATA1(19) => DATA1(19), 
                           DATA1(18) => DATA1(18), DATA1(17) => n35, DATA1(16) 
                           => DATA1(16), DATA1(15) => n48_port, DATA1(14) => 
                           n34, DATA1(13) => n60_port, DATA1(12) => DATA1(12), 
                           DATA1(11) => DATA1(11), DATA1(10) => DATA1(10), 
                           DATA1(9) => n37, DATA1(8) => n89_port, DATA1(7) => 
                           DATA1(7), DATA1(6) => n53_port, DATA1(5) => n31, 
                           DATA1(4) => DATA1(4), DATA1(3) => DATA1(3), DATA1(2)
                           => n80_port, DATA1(1) => n129, DATA1(0) => n36, 
                           DATA2(31) => DATA2(31), DATA2(30) => n63_port, 
                           DATA2(29) => DATA2(29), DATA2(28) => DATA2(28), 
                           DATA2(27) => DATA2(27), DATA2(26) => n25, DATA2(25) 
                           => DATA2(25), DATA2(24) => DATA2(24), DATA2(23) => 
                           DATA2(23), DATA2(22) => n49_port, DATA2(21) => 
                           DATA2(21), DATA2(20) => n54_port, DATA2(19) => 
                           DATA2(19), DATA2(18) => n62_port, DATA2(17) => n27, 
                           DATA2(16) => n30, DATA2(15) => DATA2(15), DATA2(14) 
                           => n29, DATA2(13) => n44, DATA2(12) => DATA2(12), 
                           DATA2(11) => n75_port, DATA2(10) => n71_port, 
                           DATA2(9) => n41, DATA2(8) => n39, DATA2(7) => 
                           DATA2(7), DATA2(6) => n45, DATA2(5) => n47_port, 
                           DATA2(4) => DATA2(4), DATA2(3) => DATA2(3), DATA2(2)
                           => n97_port, DATA2(1) => n67_port, DATA2(0) => 
                           n57_port, OUTPUT(31) => OUT_SHIFTER_31_port, 
                           OUTPUT(30) => OUT_SHIFTER_30_port, OUTPUT(29) => 
                           OUT_SHIFTER_29_port, OUTPUT(28) => 
                           OUT_SHIFTER_28_port, OUTPUT(27) => 
                           OUT_SHIFTER_27_port, OUTPUT(26) => 
                           OUT_SHIFTER_26_port, OUTPUT(25) => 
                           OUT_SHIFTER_25_port, OUTPUT(24) => 
                           OUT_SHIFTER_24_port, OUTPUT(23) => 
                           OUT_SHIFTER_23_port, OUTPUT(22) => 
                           OUT_SHIFTER_22_port, OUTPUT(21) => 
                           OUT_SHIFTER_21_port, OUTPUT(20) => 
                           OUT_SHIFTER_20_port, OUTPUT(19) => 
                           OUT_SHIFTER_19_port, OUTPUT(18) => 
                           OUT_SHIFTER_18_port, OUTPUT(17) => 
                           OUT_SHIFTER_17_port, OUTPUT(16) => 
                           OUT_SHIFTER_16_port, OUTPUT(15) => 
                           OUT_SHIFTER_15_port, OUTPUT(14) => 
                           OUT_SHIFTER_14_port, OUTPUT(13) => 
                           OUT_SHIFTER_13_port, OUTPUT(12) => 
                           OUT_SHIFTER_12_port, OUTPUT(11) => 
                           OUT_SHIFTER_11_port, OUTPUT(10) => 
                           OUT_SHIFTER_10_port, OUTPUT(9) => OUT_SHIFTER_9_port
                           , OUTPUT(8) => OUT_SHIFTER_8_port, OUTPUT(7) => 
                           OUT_SHIFTER_7_port, OUTPUT(6) => OUT_SHIFTER_6_port,
                           OUTPUT(5) => OUT_SHIFTER_5_port, OUTPUT(4) => 
                           OUT_SHIFTER_4_port, OUTPUT(3) => OUT_SHIFTER_3_port,
                           OUTPUT(2) => OUT_SHIFTER_2_port, OUTPUT(1) => 
                           OUT_SHIFTER_1_port, OUTPUT(0) => OUT_SHIFTER_0_port)
                           ;
   sub_66 : ALU_N32_DW01_sub_2 port map( A(31) => DATA1(31), A(30) => DATA1(30)
                           , A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => n26, 
                           B(7) => DATA2(7), B(6) => DATA2(6), B(5) => DATA2(5)
                           , B(4) => DATA2(4), B(3) => DATA2(3), B(2) => 
                           DATA2(2), B(1) => n43, B(0) => DATA2(0), CI => n11, 
                           DIFF(31) => N110, DIFF(30) => N109, DIFF(29) => N108
                           , DIFF(28) => N107, DIFF(27) => N106, DIFF(26) => 
                           N105, DIFF(25) => N104, DIFF(24) => N103, DIFF(23) 
                           => N102, DIFF(22) => N101, DIFF(21) => N100, 
                           DIFF(20) => N99, DIFF(19) => N98, DIFF(18) => N97, 
                           DIFF(17) => N96, DIFF(16) => N95, DIFF(15) => N94, 
                           DIFF(14) => N93, DIFF(13) => N92, DIFF(12) => N91, 
                           DIFF(11) => N90, DIFF(10) => N89, DIFF(9) => N88, 
                           DIFF(8) => N87, DIFF(7) => N86, DIFF(6) => N85, 
                           DIFF(5) => N84, DIFF(4) => N83, DIFF(3) => N82, 
                           DIFF(2) => N81, DIFF(1) => N80, DIFF(0) => N79, CO 
                           => n_1150);
   add_65 : ALU_N32_DW01_add_2 port map( A(31) => DATA1(31), A(30) => DATA1(30)
                           , A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , CI => n12, SUM(31) => N78, SUM(30) => N77, SUM(29)
                           => N76, SUM(28) => N75, SUM(27) => N74, SUM(26) => 
                           N73, SUM(25) => N72, SUM(24) => N71, SUM(23) => N70,
                           SUM(22) => N69, SUM(21) => N68, SUM(20) => N67, 
                           SUM(19) => N66, SUM(18) => N65, SUM(17) => N64, 
                           SUM(16) => N63, SUM(15) => N62, SUM(14) => N61, 
                           SUM(13) => N60, SUM(12) => N59, SUM(11) => N58, 
                           SUM(10) => N57, SUM(9) => N56, SUM(8) => N55, SUM(7)
                           => N54, SUM(6) => N53, SUM(5) => N52, SUM(4) => N51,
                           SUM(3) => N50, SUM(2) => N49, SUM(1) => N48, SUM(0) 
                           => N47, CO => n_1151);
   r59 : ALU_N32_DW01_cmp6_2 port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => n32, A(12) => DATA1(12)
                           , A(11) => DATA1(11), A(10) => DATA1(10), A(9) => 
                           n37, A(8) => n89_port, A(7) => DATA1(7), A(6) => 
                           n87_port, A(5) => n31, A(4) => n130, A(3) => 
                           n52_port, A(2) => n100_port, A(1) => n129, A(0) => 
                           n36, B(31) => DATA2(31), B(30) => DATA2(30), B(29) 
                           => DATA2(29), B(28) => DATA2(28), B(27) => DATA2(27)
                           , B(26) => DATA2(26), B(25) => DATA2(25), B(24) => 
                           DATA2(24), B(23) => DATA2(23), B(22) => DATA2(22), 
                           B(21) => DATA2(21), B(20) => DATA2(20), B(19) => 
                           DATA2(19), B(18) => DATA2(18), B(17) => DATA2(17), 
                           B(16) => DATA2(16), B(15) => n24, B(14) => DATA2(14)
                           , B(13) => n28, B(12) => DATA2(12), B(11) => 
                           DATA2(11), B(10) => DATA2(10), B(9) => DATA2(9), 
                           B(8) => n46, B(7) => DATA2(7), B(6) => n45, B(5) => 
                           DATA2(5), B(4) => n68_port, B(3) => n50_port, B(2) 
                           => n112_port, B(1) => n67_port, B(0) => n57_port, TC
                           => n13, LT => n_1152, GT => n_1153, EQ => n_1154, LE
                           => N111, GE => N112, NE => n_1155);
   ne_72 : ALU_N32_DW01_cmp6_3 port map( A(31) => DATA1(31), A(30) => DATA1(30)
                           , A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => n38, A(18) => DATA1(18), A(17) => n61_port,
                           A(16) => n20, A(15) => n48_port, A(14) => n76_port, 
                           A(13) => n60_port, A(12) => n51_port, A(11) => 
                           DATA1(11), A(10) => DATA1(10), A(9) => n98_port, 
                           A(8) => n113_port, A(7) => n55_port, A(6) => 
                           n74_port, A(5) => n69_port, A(4) => n1, A(3) => 
                           n52_port, A(2) => n100_port, A(1) => n129, A(0) => 
                           n36, B(31) => DATA2(31), B(30) => DATA2(30), B(29) 
                           => DATA2(29), B(28) => DATA2(28), B(27) => DATA2(27)
                           , B(26) => DATA2(26), B(25) => DATA2(25), B(24) => 
                           DATA2(24), B(23) => DATA2(23), B(22) => DATA2(22), 
                           B(21) => DATA2(21), B(20) => DATA2(20), B(19) => 
                           DATA2(19), B(18) => DATA2(18), B(17) => n27, B(16) 
                           => n30, B(15) => DATA2(15), B(14) => n29, B(13) => 
                           n44, B(12) => DATA2(12), B(11) => DATA2(11), B(10) 
                           => DATA2(10), B(9) => n41, B(8) => n39, B(7) => 
                           DATA2(7), B(6) => n45, B(5) => n47_port, B(4) => 
                           n99_port, B(3) => n65_port, B(2) => n112_port, B(1) 
                           => n85_port, B(0) => n57_port, TC => n10, LT => 
                           n_1156, GT => n_1157, EQ => n_1158, LE => n_1159, GE
                           => n_1160, NE => N113);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26 is

   port( NOT_EXT_IMM : in std_logic_vector (25 downto 0);  SIGNED_IMM, IS_JUMP 
         : in std_logic;  EXT_IMM : out std_logic_vector (31 downto 0));

end EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26;

architecture SYN_BEHAVIOR of EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal EXT_IMM_31_port, EXT_IMM_25_port, EXT_IMM_24_port, EXT_IMM_23_port, 
      EXT_IMM_22_port, EXT_IMM_21_port, EXT_IMM_20_port, EXT_IMM_19_port, 
      EXT_IMM_18_port, EXT_IMM_17_port, EXT_IMM_16_port, n3, n4, n5, n6, n7, n8
      , n9, n10, n11, n12, n13, n1, n2 : std_logic;

begin
   EXT_IMM <= ( EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, 
      EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_25_port, 
      EXT_IMM_24_port, EXT_IMM_23_port, EXT_IMM_22_port, EXT_IMM_21_port, 
      EXT_IMM_20_port, EXT_IMM_19_port, EXT_IMM_18_port, EXT_IMM_17_port, 
      EXT_IMM_16_port, NOT_EXT_IMM(15), NOT_EXT_IMM(14), NOT_EXT_IMM(13), 
      NOT_EXT_IMM(12), NOT_EXT_IMM(11), NOT_EXT_IMM(10), NOT_EXT_IMM(9), 
      NOT_EXT_IMM(8), NOT_EXT_IMM(7), NOT_EXT_IMM(6), NOT_EXT_IMM(5), 
      NOT_EXT_IMM(4), NOT_EXT_IMM(3), NOT_EXT_IMM(2), NOT_EXT_IMM(1), 
      NOT_EXT_IMM(0) );
   
   U24 : NAND3_X1 port map( A1 => NOT_EXT_IMM(25), A2 => IS_JUMP, A3 => 
                           SIGNED_IMM, ZN => n4);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n6, ZN => EXT_IMM_23_port);
   U3 : NAND2_X1 port map( A1 => NOT_EXT_IMM(23), A2 => IS_JUMP, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n5, ZN => EXT_IMM_24_port);
   U5 : NAND2_X1 port map( A1 => NOT_EXT_IMM(24), A2 => IS_JUMP, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n8, ZN => EXT_IMM_21_port);
   U7 : NAND2_X1 port map( A1 => NOT_EXT_IMM(21), A2 => IS_JUMP, ZN => n8);
   U8 : NAND2_X1 port map( A1 => n3, A2 => n10, ZN => EXT_IMM_19_port);
   U9 : NAND2_X1 port map( A1 => NOT_EXT_IMM(19), A2 => IS_JUMP, ZN => n10);
   U10 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n3, ZN => EXT_IMM_25_port)
                           ;
   U11 : INV_X1 port map( A => NOT_EXT_IMM(25), ZN => n1);
   U12 : NAND2_X1 port map( A1 => n3, A2 => n12, ZN => EXT_IMM_17_port);
   U13 : NAND2_X1 port map( A1 => NOT_EXT_IMM(17), A2 => IS_JUMP, ZN => n12);
   U14 : NAND2_X1 port map( A1 => n3, A2 => n11, ZN => EXT_IMM_18_port);
   U15 : NAND2_X1 port map( A1 => NOT_EXT_IMM(18), A2 => IS_JUMP, ZN => n11);
   U16 : NAND2_X1 port map( A1 => n3, A2 => n13, ZN => EXT_IMM_16_port);
   U17 : NAND2_X1 port map( A1 => NOT_EXT_IMM(16), A2 => IS_JUMP, ZN => n13);
   U18 : NAND2_X1 port map( A1 => n3, A2 => n7, ZN => EXT_IMM_22_port);
   U19 : NAND2_X1 port map( A1 => NOT_EXT_IMM(22), A2 => IS_JUMP, ZN => n7);
   U20 : NAND2_X1 port map( A1 => n3, A2 => n9, ZN => EXT_IMM_20_port);
   U21 : NAND2_X1 port map( A1 => NOT_EXT_IMM(20), A2 => IS_JUMP, ZN => n9);
   U22 : NAND3_X1 port map( A1 => SIGNED_IMM, A2 => n2, A3 => NOT_EXT_IMM(15), 
                           ZN => n3);
   U23 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => EXT_IMM_31_port);
   U25 : INV_X1 port map( A => IS_JUMP, ZN => n2);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REGISTER_FILE_NBIT32_NREG32 is

   port( CLK, RST, EN, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 :
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0));

end REGISTER_FILE_NBIT32_NREG32;

architecture SYN_BEHAVIOR of REGISTER_FILE_NBIT32_NREG32 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
      n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
      n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
      n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, 
      n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
      n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
      n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, 
      n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
      n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
      n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
      n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
      n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, 
      n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
      n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
      n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
      n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, 
      n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
      n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, 
      n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, 
      n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
      n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
      n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, 
      n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, 
      n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
      n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, 
      n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, 
      n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, 
      n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
      n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, 
      n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
      n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, 
      n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
      n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, 
      n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
      n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, 
      n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, 
      n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, 
      n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, 
      n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, 
      n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, 
      n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, 
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, 
      n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
      n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, 
      n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, 
      n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, 
      n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, 
      n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, 
      n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, 
      n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, 
      n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, 
      n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, 
      n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, 
      n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, 
      n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, 
      n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, 
      n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, 
      n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, 
      n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, 
      n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, 
      n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, 
      n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, 
      n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, 
      n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, 
      n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, 
      n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, 
      n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, 
      n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, 
      n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, 
      n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, 
      n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, 
      n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, 
      n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, 
      n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, 
      n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, 
      n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, 
      n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, 
      n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, 
      n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, 
      n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, 
      n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, 
      n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
      n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
      n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
      n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, 
      n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, 
      n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
      n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, 
      n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
      n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, 
      n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
      n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, 
      n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, 
      n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, 
      n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, 
      n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
      n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
      n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, 
      n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, 
      n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, 
      n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, 
      n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
      n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, 
      n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, 
      n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, 
      n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, 
      n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, 
      n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, 
      n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, 
      n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, 
      n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, 
      n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, 
      n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, 
      n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, 
      n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, 
      n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, 
      n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, 
      n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, 
      n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, 
      n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, 
      n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, 
      n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, 
      n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, 
      n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, 
      n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, 
      n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, 
      n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, 
      n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, 
      n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, 
      n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, 
      n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, 
      n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, 
      n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, 
      n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, 
      n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, 
      n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, 
      n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, 
      n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, 
      n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, 
      n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, 
      n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, 
      n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
      n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
      n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, 
      n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, 
      n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, 
      n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, 
      n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, 
      n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, 
      n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, 
      n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, 
      n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, 
      n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, 
      n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, 
      n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, 
      n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, 
      n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, 
      n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, 
      n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, 
      n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
      n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, 
      n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
      n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, 
      n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, 
      n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, 
      n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, 
      n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, 
      n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, 
      n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, 
      n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
      n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, 
      n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
      n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, 
      n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, 
      n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, 
      n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, 
      n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, 
      n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, 
      n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, 
      n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, 
      n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, 
      n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
      n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, 
      n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, 
      n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, 
      n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, 
      n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, 
      n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, 
      n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, 
      n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, 
      n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, 
      n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, 
      n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, 
      n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, 
      n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, 
      n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, 
      n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, 
      n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, 
      n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, 
      n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, 
      n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, 
      n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
      n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, 
      n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, 
      n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, 
      n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, 
      n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, 
      n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, 
      n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, 
      n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, 
      n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, 
      n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, 
      n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, 
      n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, 
      n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, 
      n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, 
      n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, 
      n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, 
      n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, 
      n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, 
      n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, 
      n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
      n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, 
      n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, 
      n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
      n2525, n2526, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, 
      n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, 
      n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, 
      n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
      n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, 
      n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
      n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
      n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
      n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
      n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, 
      n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
      n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
      n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
      n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, 
      n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
      n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, 
      n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
      n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
      n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
      n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, 
      n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
      n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
      n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, 
      n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
      n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
      n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, 
      n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, 
      n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
      n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
      n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
      n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, 
      n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, 
      n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, 
      n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
      n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
      n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, 
      n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, 
      n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, 
      n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, 
      n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, 
      n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, 
      n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, 
      n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, 
      n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, 
      n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, 
      n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, 
      n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, 
      n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, 
      n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, 
      n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, 
      n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, 
      n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, 
      n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, 
      n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, 
      n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, 
      n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, 
      n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, 
      n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, 
      n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, 
      n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, 
      n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, 
      n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, 
      n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, 
      n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, 
      n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, 
      n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, 
      n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, 
      n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, 
      n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, 
      n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, 
      n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, 
      n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, 
      n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, 
      n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, 
      n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, 
      n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, 
      n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, 
      n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, 
      n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, 
      n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, 
      n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, 
      n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, 
      n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, 
      n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, 
      n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, 
      n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, 
      n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, 
      n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, 
      n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, 
      n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, 
      n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, 
      n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, 
      n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, 
      n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, 
      n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, 
      n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, 
      n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, 
      n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, 
      n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, 
      n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, 
      n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, 
      n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, 
      n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, 
      n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, 
      n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, 
      n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, 
      n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, 
      n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, 
      n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, 
      n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, 
      n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, 
      n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, 
      n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, 
      n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, 
      n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, 
      n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, 
      n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, 
      n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, 
      n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, 
      n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, 
      n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, 
      n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, 
      n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, 
      n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, 
      n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, 
      n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, 
      n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, 
      n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, 
      n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, 
      n_2180, n_2181, n_2182, n_2183, n_2184 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n3614, CK => CLK, Q => 
                           n_1161, QN => n2166);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => 
                           n_1162, QN => n2124);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => 
                           n_1163, QN => n2088);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => 
                           n_1164, QN => n2052);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => 
                           n_1165, QN => n2016);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => 
                           n_1166, QN => n1981);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => 
                           n_1167, QN => n1946);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => 
                           n_1168, QN => n1910);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => 
                           n_1169, QN => n1874);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => 
                           n_1170, QN => n1838);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => 
                           n_1171, QN => n1802);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => 
                           n_1172, QN => n1766);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => 
                           n_1173, QN => n1730);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => 
                           n_1174, QN => n1695);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => 
                           n_1175, QN => n1659);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => 
                           n_1176, QN => n1623);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => 
                           n_1177, QN => n1588);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => 
                           n_1178, QN => n1553);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => 
                           n_1179, QN => n1517);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => 
                           n_1180, QN => n1482);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => 
                           n_1181, QN => n1447);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => 
                           n_1182, QN => n1412);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => n_1183
                           , QN => n1377);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => n_1184
                           , QN => n1342);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => n_1185
                           , QN => n1306);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => n_1186
                           , QN => n1270);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => n_1187
                           , QN => n1234);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => n_1188
                           , QN => n1198);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => n_1189
                           , QN => n1162);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => n_1190
                           , QN => n1126);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => n_1191
                           , QN => n1090);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => n_1192
                           , QN => n1052);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => 
                           n_1193, QN => n2168);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => 
                           n_1194, QN => n2125);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => 
                           n_1195, QN => n2089);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => 
                           n_1196, QN => n2053);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => 
                           n_1197, QN => n2017);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => 
                           n_1198, QN => n1982);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => 
                           n_1199, QN => n1947);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => 
                           n_1200, QN => n1911);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => 
                           n_1201, QN => n1875);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => 
                           n_1202, QN => n1839);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => 
                           n_1203, QN => n1803);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => 
                           n_1204, QN => n1767);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => 
                           n_1205, QN => n1731);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => 
                           n_1206, QN => n1696);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => 
                           n_1207, QN => n1660);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => 
                           n_1208, QN => n1624);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => 
                           n_1209, QN => n1589);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => 
                           n_1210, QN => n1554);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => 
                           n_1211, QN => n1518);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => 
                           n_1212, QN => n1483);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => 
                           n_1213, QN => n1448);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => 
                           n_1214, QN => n1413);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => n_1215
                           , QN => n1378);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => n_1216
                           , QN => n1343);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => n_1217
                           , QN => n1307);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => n_1218
                           , QN => n1271);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => n_1219
                           , QN => n1235);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => n_1220
                           , QN => n1199);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => n_1221
                           , QN => n1163);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => n_1222
                           , QN => n1127);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => n_1223
                           , QN => n1091);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => n_1224
                           , QN => n1053);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => n4356
                           , QN => n_1225);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => n4353
                           , QN => n_1226);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => n4351
                           , QN => n_1227);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => n4349
                           , QN => n_1228);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => n4347
                           , QN => n_1229);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => n4345
                           , QN => n_1230);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => n4343
                           , QN => n_1231);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => n4341
                           , QN => n_1232);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => n4339
                           , QN => n_1233);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => n4337
                           , QN => n_1234);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => n4335
                           , QN => n_1235);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => n4333
                           , QN => n_1236);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => n4331
                           , QN => n_1237);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => n4329
                           , QN => n_1238);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => n4327
                           , QN => n_1239);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => n4325
                           , QN => n_1240);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => n4323
                           , QN => n_1241);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => n4321
                           , QN => n_1242);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => n4319
                           , QN => n_1243);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => n4317
                           , QN => n_1244);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => n4315
                           , QN => n_1245);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => n4313
                           , QN => n_1246);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => n4311,
                           QN => n_1247);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => n4309,
                           QN => n_1248);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n3526, CK => CLK, Q => n4307,
                           QN => n_1249);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => n4305,
                           QN => n_1250);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => n4303,
                           QN => n_1251);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => n4301,
                           QN => n_1252);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => n4299,
                           QN => n_1253);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => n4297,
                           QN => n_1254);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => n4295,
                           QN => n_1255);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => n4293,
                           QN => n_1256);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => n4290
                           , QN => n_1257);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => n4288
                           , QN => n_1258);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => n4287
                           , QN => n_1259);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => n4286
                           , QN => n_1260);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => n4285
                           , QN => n_1261);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => n4284
                           , QN => n_1262);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => n4283
                           , QN => n_1263);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => n4282
                           , QN => n_1264);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => n4281
                           , QN => n_1265);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => n4280
                           , QN => n_1266);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => n4279
                           , QN => n_1267);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => n4278
                           , QN => n_1268);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => n4277
                           , QN => n_1269);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => n4276
                           , QN => n_1270);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => n4275
                           , QN => n_1271);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => n4274
                           , QN => n_1272);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => n4273
                           , QN => n_1273);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => n4272
                           , QN => n_1274);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => n4271
                           , QN => n_1275);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => n4270
                           , QN => n_1276);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => n4269
                           , QN => n_1277);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => n4268
                           , QN => n_1278);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => n4267,
                           QN => n_1279);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => n4266,
                           QN => n_1280);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => n4265,
                           QN => n_1281);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => n4264,
                           QN => n_1282);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => n4263,
                           QN => n_1283);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => n4262,
                           QN => n_1284);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => n4261,
                           QN => n_1285);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => n4260,
                           QN => n_1286);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => n4259,
                           QN => n_1287);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => n4258,
                           QN => n_1288);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => 
                           n_1289, QN => n2161);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => 
                           n_1290, QN => n2121);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => 
                           n_1291, QN => n2085);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => 
                           n_1292, QN => n2049);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => 
                           n_1293, QN => n2013);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => 
                           n_1294, QN => n1978);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => 
                           n_1295, QN => n1943);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => 
                           n_1296, QN => n1907);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => 
                           n_1297, QN => n1871);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => 
                           n_1298, QN => n1835);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => 
                           n_1299, QN => n1799);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => 
                           n_1300, QN => n1763);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => 
                           n_1301, QN => n1727);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => 
                           n_1302, QN => n1692);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n3472, CK => CLK, Q => 
                           n_1303, QN => n1656);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => 
                           n_1304, QN => n1620);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => 
                           n_1305, QN => n1585);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => 
                           n_1306, QN => n1550);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => 
                           n_1307, QN => n1514);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => 
                           n_1308, QN => n1479);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => 
                           n_1309, QN => n1444);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => 
                           n_1310, QN => n1409);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => n_1311
                           , QN => n1374);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => n_1312
                           , QN => n1339);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => n_1313
                           , QN => n1303);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => n_1314
                           , QN => n1267);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => n_1315
                           , QN => n1231);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => n_1316
                           , QN => n1195);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => n_1317
                           , QN => n1159);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => n_1318
                           , QN => n1123);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => n_1319
                           , QN => n1087);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => n_1320
                           , QN => n1049);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => 
                           n_1321, QN => n2163);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => 
                           n_1322, QN => n2122);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => 
                           n_1323, QN => n2086);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => 
                           n_1324, QN => n2050);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => 
                           n_1325, QN => n2014);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => 
                           n_1326, QN => n1979);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => 
                           n_1327, QN => n1944);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => 
                           n_1328, QN => n1908);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => 
                           n_1329, QN => n1872);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => 
                           n_1330, QN => n1836);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => 
                           n_1331, QN => n1800);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => 
                           n_1332, QN => n1764);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => 
                           n_1333, QN => n1728);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => 
                           n_1334, QN => n1693);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => 
                           n_1335, QN => n1657);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => 
                           n_1336, QN => n1621);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => 
                           n_1337, QN => n1586);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => 
                           n_1338, QN => n1551);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => 
                           n_1339, QN => n1515);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => 
                           n_1340, QN => n1480);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => 
                           n_1341, QN => n1445);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => 
                           n_1342, QN => n1410);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => n_1343
                           , QN => n1375);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => n_1344
                           , QN => n1340);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => n_1345
                           , QN => n1304);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => n_1346
                           , QN => n1268);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => n_1347
                           , QN => n1232);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => n_1348
                           , QN => n1196);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => n_1349
                           , QN => n1160);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => n_1350
                           , QN => n1124);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => n_1351
                           , QN => n1088);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => n_1352
                           , QN => n1050);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => n4185
                           , QN => n_1353);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => n4183
                           , QN => n_1354);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => n4182
                           , QN => n_1355);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => n4181
                           , QN => n_1356);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => n4180
                           , QN => n_1357);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => n4179
                           , QN => n_1358);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => n4178
                           , QN => n_1359);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => n4177
                           , QN => n_1360);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => n4176
                           , QN => n_1361);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => n4175
                           , QN => n_1362);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => n4174
                           , QN => n_1363);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => n4173
                           , QN => n_1364);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => n4172
                           , QN => n_1365);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => n4171
                           , QN => n_1366);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => n4170
                           , QN => n_1367);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => n4169
                           , QN => n_1368);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => n4168
                           , QN => n_1369);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => n4167
                           , QN => n_1370);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => n4166
                           , QN => n_1371);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => n4165
                           , QN => n_1372);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => n4164
                           , QN => n_1373);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => n4163
                           , QN => n_1374);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => n4162,
                           QN => n_1375);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => n4161,
                           QN => n_1376);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => n4160,
                           QN => n_1377);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => n4159,
                           QN => n_1378);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => n4158,
                           QN => n_1379);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => n4157,
                           QN => n_1380);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => n4156,
                           QN => n_1381);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => n4155,
                           QN => n_1382);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => n4154,
                           QN => n_1383);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => n4153,
                           QN => n_1384);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => n4150
                           , QN => n_1385);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => n4148
                           , QN => n_1386);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => n4147
                           , QN => n_1387);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => n4146
                           , QN => n_1388);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => n4145
                           , QN => n_1389);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => n4144
                           , QN => n_1390);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => n4143
                           , QN => n_1391);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => n4142
                           , QN => n_1392);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => n4141
                           , QN => n_1393);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => n4140
                           , QN => n_1394);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => n4139
                           , QN => n_1395);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => n4138
                           , QN => n_1396);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => n4137
                           , QN => n_1397);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => n4136
                           , QN => n_1398);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => n4135
                           , QN => n_1399);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => n4134
                           , QN => n_1400);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => n4133
                           , QN => n_1401);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => n4132
                           , QN => n_1402);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => n4131
                           , QN => n_1403);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => n4130
                           , QN => n_1404);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => n4129
                           , QN => n_1405);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => n4128
                           , QN => n_1406);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => n4127,
                           QN => n_1407);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => n4126,
                           QN => n_1408);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => n4125,
                           QN => n_1409);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => n4124,
                           QN => n_1410);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => n4123,
                           QN => n_1411);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => n4122,
                           QN => n_1412);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => n4121,
                           QN => n_1413);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => n4120,
                           QN => n_1414);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => n4119,
                           QN => n_1415);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => n4118,
                           QN => n_1416);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => 
                           n_1417, QN => n2156);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => 
                           n_1418, QN => n2118);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => 
                           n_1419, QN => n2082);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => 
                           n_1420, QN => n2046);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => 
                           n_1421, QN => n2010);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => 
                           n_1422, QN => n1975);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => 
                           n_1423, QN => n1940);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => 
                           n_1424, QN => n1904);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => 
                           n_1425, QN => n1868);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => 
                           n_1426, QN => n1832);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => 
                           n_1427, QN => n1796);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => 
                           n_1428, QN => n1760);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => 
                           n_1429, QN => n1724);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => 
                           n_1430, QN => n1689);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => 
                           n_1431, QN => n1653);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => 
                           n_1432, QN => n1617);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => 
                           n_1433, QN => n1582);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => 
                           n_1434, QN => n1547);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => 
                           n_1435, QN => n1511);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => 
                           n_1436, QN => n1476);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => 
                           n_1437, QN => n1441);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => 
                           n_1438, QN => n1406);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => n_1439
                           , QN => n1371);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => n_1440
                           , QN => n1336);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => n_1441
                           , QN => n1300);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => n_1442
                           , QN => n1264);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => n_1443
                           , QN => n1228);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => n_1444
                           , QN => n1192);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => n_1445
                           , QN => n1156);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => n_1446
                           , QN => n1120);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => n_1447
                           , QN => n1084);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => n_1448
                           , QN => n1045);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3326, CK => CLK, Q => 
                           n_1449, QN => n2158);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => 
                           n_1450, QN => n2119);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => 
                           n_1451, QN => n2083);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => 
                           n_1452, QN => n2047);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => 
                           n_1453, QN => n2011);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => 
                           n_1454, QN => n1976);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => 
                           n_1455, QN => n1941);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => 
                           n_1456, QN => n1905);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => 
                           n_1457, QN => n1869);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => 
                           n_1458, QN => n1833);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => 
                           n_1459, QN => n1797);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => 
                           n_1460, QN => n1761);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => 
                           n_1461, QN => n1725);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => 
                           n_1462, QN => n1690);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => 
                           n_1463, QN => n1654);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => 
                           n_1464, QN => n1618);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => 
                           n_1465, QN => n1583);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => 
                           n_1466, QN => n1548);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => 
                           n_1467, QN => n1512);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => 
                           n_1468, QN => n1477);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => 
                           n_1469, QN => n1442);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => 
                           n_1470, QN => n1407);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => n_1471
                           , QN => n1372);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => n_1472
                           , QN => n1337);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => n_1473
                           , QN => n1301);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => n_1474
                           , QN => n1265);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => n_1475
                           , QN => n1229);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => n_1476
                           , QN => n1193);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => n_1477
                           , QN => n1157);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => n_1478
                           , QN => n1121);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => n_1479
                           , QN => n1085);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => n_1480
                           , QN => n1046);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => 
                           n4044, QN => n_1481);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => 
                           n4042, QN => n_1482);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => 
                           n4041, QN => n_1483);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => 
                           n4040, QN => n_1484);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => 
                           n4039, QN => n_1485);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3289, CK => CLK, Q => 
                           n4038, QN => n_1486);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => 
                           n4037, QN => n_1487);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => 
                           n4036, QN => n_1488);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => 
                           n4035, QN => n_1489);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => 
                           n4034, QN => n_1490);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => 
                           n4033, QN => n_1491);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => 
                           n4032, QN => n_1492);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => 
                           n4031, QN => n_1493);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => 
                           n4030, QN => n_1494);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => 
                           n4029, QN => n_1495);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => 
                           n4028, QN => n_1496);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => 
                           n4027, QN => n_1497);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => 
                           n4026, QN => n_1498);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => 
                           n4025, QN => n_1499);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => 
                           n4024, QN => n_1500);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3274, CK => CLK, Q => 
                           n4023, QN => n_1501);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3273, CK => CLK, Q => 
                           n4022, QN => n_1502);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3272, CK => CLK, Q => n4021
                           , QN => n_1503);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3271, CK => CLK, Q => n4020
                           , QN => n_1504);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3270, CK => CLK, Q => n4019
                           , QN => n_1505);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3269, CK => CLK, Q => n4018
                           , QN => n_1506);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3268, CK => CLK, Q => n4017
                           , QN => n_1507);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3267, CK => CLK, Q => n4016
                           , QN => n_1508);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3266, CK => CLK, Q => n4015
                           , QN => n_1509);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3265, CK => CLK, Q => n4014
                           , QN => n_1510);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3264, CK => CLK, Q => n4013
                           , QN => n_1511);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3263, CK => CLK, Q => n4012
                           , QN => n_1512);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3262, CK => CLK, Q => 
                           n4010, QN => n_1513);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => 
                           n4008, QN => n_1514);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => 
                           n4007, QN => n_1515);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => 
                           n4006, QN => n_1516);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => 
                           n4005, QN => n_1517);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => 
                           n4004, QN => n_1518);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => 
                           n4003, QN => n_1519);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => 
                           n4002, QN => n_1520);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => 
                           n4001, QN => n_1521);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => 
                           n4000, QN => n_1522);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => 
                           n3999, QN => n_1523);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => 
                           n3998, QN => n_1524);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => 
                           n3997, QN => n_1525);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => 
                           n3996, QN => n_1526);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => 
                           n3995, QN => n_1527);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => 
                           n3994, QN => n_1528);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => 
                           n3993, QN => n_1529);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => 
                           n3992, QN => n_1530);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => 
                           n3991, QN => n_1531);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => 
                           n3990, QN => n_1532);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => 
                           n3989, QN => n_1533);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => 
                           n3988, QN => n_1534);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => n3987
                           , QN => n_1535);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => n3986
                           , QN => n_1536);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => n3985
                           , QN => n_1537);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => n3984
                           , QN => n_1538);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => n3983
                           , QN => n_1539);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => n3982
                           , QN => n_1540);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => n3981
                           , QN => n_1541);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => n3980
                           , QN => n_1542);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => n3979
                           , QN => n_1543);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => n3978
                           , QN => n_1544);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => 
                           n_1545, QN => n2151);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => 
                           n_1546, QN => n2115);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => 
                           n_1547, QN => n2079);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => 
                           n_1548, QN => n2043);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => 
                           n_1549, QN => n2007);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => 
                           n_1550, QN => n1972);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => 
                           n_1551, QN => n1937);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => 
                           n_1552, QN => n1901);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => 
                           n_1553, QN => n1865);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => 
                           n_1554, QN => n1829);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => 
                           n_1555, QN => n1793);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => 
                           n_1556, QN => n1757);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => 
                           n_1557, QN => n1721);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => 
                           n_1558, QN => n1686);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => 
                           n_1559, QN => n1650);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => 
                           n_1560, QN => n1614);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => 
                           n_1561, QN => n1579);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => 
                           n_1562, QN => n1544);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => 
                           n_1563, QN => n1508);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => 
                           n_1564, QN => n1473);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => 
                           n_1565, QN => n1438);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => 
                           n_1566, QN => n1403);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3208, CK => CLK, Q => 
                           n_1567, QN => n1368);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => 
                           n_1568, QN => n1333);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => 
                           n_1569, QN => n1297);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => 
                           n_1570, QN => n1261);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => 
                           n_1571, QN => n1225);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => 
                           n_1572, QN => n1189);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => 
                           n_1573, QN => n1153);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => 
                           n_1574, QN => n1117);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => 
                           n_1575, QN => n1081);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => 
                           n_1576, QN => n1040);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => 
                           n_1577, QN => n2153);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => 
                           n_1578, QN => n2116);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => 
                           n_1579, QN => n2080);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3195, CK => CLK, Q => 
                           n_1580, QN => n2044);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3194, CK => CLK, Q => 
                           n_1581, QN => n2008);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3193, CK => CLK, Q => 
                           n_1582, QN => n1973);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3192, CK => CLK, Q => 
                           n_1583, QN => n1938);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3191, CK => CLK, Q => 
                           n_1584, QN => n1902);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3190, CK => CLK, Q => 
                           n_1585, QN => n1866);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3189, CK => CLK, Q => 
                           n_1586, QN => n1830);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3188, CK => CLK, Q => 
                           n_1587, QN => n1794);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3187, CK => CLK, Q => 
                           n_1588, QN => n1758);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3186, CK => CLK, Q => 
                           n_1589, QN => n1722);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3185, CK => CLK, Q => 
                           n_1590, QN => n1687);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3184, CK => CLK, Q => 
                           n_1591, QN => n1651);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3183, CK => CLK, Q => 
                           n_1592, QN => n1615);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3182, CK => CLK, Q => 
                           n_1593, QN => n1580);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3181, CK => CLK, Q => 
                           n_1594, QN => n1545);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3180, CK => CLK, Q => 
                           n_1595, QN => n1509);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3179, CK => CLK, Q => 
                           n_1596, QN => n1474);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3178, CK => CLK, Q => 
                           n_1597, QN => n1439);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3177, CK => CLK, Q => 
                           n_1598, QN => n1404);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3176, CK => CLK, Q => 
                           n_1599, QN => n1369);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3175, CK => CLK, Q => 
                           n_1600, QN => n1334);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3174, CK => CLK, Q => 
                           n_1601, QN => n1298);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3173, CK => CLK, Q => 
                           n_1602, QN => n1262);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3172, CK => CLK, Q => 
                           n_1603, QN => n1226);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3171, CK => CLK, Q => 
                           n_1604, QN => n1190);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3170, CK => CLK, Q => 
                           n_1605, QN => n1154);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3169, CK => CLK, Q => 
                           n_1606, QN => n1118);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3168, CK => CLK, Q => 
                           n_1607, QN => n1082);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3167, CK => CLK, Q => 
                           n_1608, QN => n1041);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3166, CK => CLK, Q => 
                           n3908, QN => n_1609);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3165, CK => CLK, Q => 
                           n3906, QN => n_1610);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3164, CK => CLK, Q => 
                           n3905, QN => n_1611);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3163, CK => CLK, Q => 
                           n3904, QN => n_1612);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3162, CK => CLK, Q => 
                           n3903, QN => n_1613);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3161, CK => CLK, Q => 
                           n3902, QN => n_1614);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3160, CK => CLK, Q => 
                           n3901, QN => n_1615);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3159, CK => CLK, Q => 
                           n3900, QN => n_1616);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3158, CK => CLK, Q => 
                           n3899, QN => n_1617);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3157, CK => CLK, Q => 
                           n3898, QN => n_1618);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3156, CK => CLK, Q => 
                           n3897, QN => n_1619);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3155, CK => CLK, Q => 
                           n3896, QN => n_1620);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3154, CK => CLK, Q => 
                           n3895, QN => n_1621);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3153, CK => CLK, Q => 
                           n3894, QN => n_1622);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3152, CK => CLK, Q => 
                           n3893, QN => n_1623);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3151, CK => CLK, Q => 
                           n3892, QN => n_1624);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3150, CK => CLK, Q => 
                           n3891, QN => n_1625);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3149, CK => CLK, Q => 
                           n3890, QN => n_1626);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3148, CK => CLK, Q => 
                           n3889, QN => n_1627);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3147, CK => CLK, Q => 
                           n3888, QN => n_1628);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3146, CK => CLK, Q => 
                           n3887, QN => n_1629);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3145, CK => CLK, Q => 
                           n3886, QN => n_1630);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3144, CK => CLK, Q => n3885
                           , QN => n_1631);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3143, CK => CLK, Q => n3884
                           , QN => n_1632);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3142, CK => CLK, Q => n3883
                           , QN => n_1633);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3141, CK => CLK, Q => n3882
                           , QN => n_1634);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3140, CK => CLK, Q => n3881
                           , QN => n_1635);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3139, CK => CLK, Q => n3880
                           , QN => n_1636);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3138, CK => CLK, Q => n3879
                           , QN => n_1637);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3137, CK => CLK, Q => n3878
                           , QN => n_1638);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3136, CK => CLK, Q => n3877
                           , QN => n_1639);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3135, CK => CLK, Q => n3876
                           , QN => n_1640);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3134, CK => CLK, Q => 
                           n3874, QN => n_1641);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3133, CK => CLK, Q => 
                           n3872, QN => n_1642);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3132, CK => CLK, Q => 
                           n3871, QN => n_1643);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3131, CK => CLK, Q => 
                           n3870, QN => n_1644);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3130, CK => CLK, Q => 
                           n3869, QN => n_1645);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3129, CK => CLK, Q => 
                           n3868, QN => n_1646);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3128, CK => CLK, Q => 
                           n3867, QN => n_1647);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3127, CK => CLK, Q => 
                           n3866, QN => n_1648);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3126, CK => CLK, Q => 
                           n3865, QN => n_1649);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3125, CK => CLK, Q => 
                           n3864, QN => n_1650);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3124, CK => CLK, Q => 
                           n3863, QN => n_1651);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3123, CK => CLK, Q => 
                           n3862, QN => n_1652);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3122, CK => CLK, Q => 
                           n3861, QN => n_1653);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3121, CK => CLK, Q => 
                           n3860, QN => n_1654);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3120, CK => CLK, Q => 
                           n3859, QN => n_1655);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3119, CK => CLK, Q => 
                           n3858, QN => n_1656);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3118, CK => CLK, Q => 
                           n3857, QN => n_1657);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3117, CK => CLK, Q => 
                           n3856, QN => n_1658);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3116, CK => CLK, Q => 
                           n3855, QN => n_1659);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3115, CK => CLK, Q => 
                           n3854, QN => n_1660);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3114, CK => CLK, Q => 
                           n3853, QN => n_1661);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3113, CK => CLK, Q => 
                           n3852, QN => n_1662);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3112, CK => CLK, Q => n3851
                           , QN => n_1663);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3111, CK => CLK, Q => n3850
                           , QN => n_1664);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3110, CK => CLK, Q => n3849
                           , QN => n_1665);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3109, CK => CLK, Q => n3848
                           , QN => n_1666);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3108, CK => CLK, Q => n3847
                           , QN => n_1667);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3107, CK => CLK, Q => n3846
                           , QN => n_1668);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3106, CK => CLK, Q => n3845
                           , QN => n_1669);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3105, CK => CLK, Q => n3844
                           , QN => n_1670);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3104, CK => CLK, Q => n3843
                           , QN => n_1671);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3103, CK => CLK, Q => n3842
                           , QN => n_1672);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3102, CK => CLK, Q => 
                           n_1673, QN => n2190);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3101, CK => CLK, Q => 
                           n_1674, QN => n2140);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3100, CK => CLK, Q => 
                           n_1675, QN => n2104);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3099, CK => CLK, Q => 
                           n_1676, QN => n2068);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3098, CK => CLK, Q => 
                           n_1677, QN => n2032);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3097, CK => CLK, Q => 
                           n_1678, QN => n1997);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3096, CK => CLK, Q => 
                           n_1679, QN => n1962);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3095, CK => CLK, Q => 
                           n_1680, QN => n1926);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3094, CK => CLK, Q => 
                           n_1681, QN => n1890);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3093, CK => CLK, Q => 
                           n_1682, QN => n1854);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3092, CK => CLK, Q => 
                           n_1683, QN => n1818);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3091, CK => CLK, Q => 
                           n_1684, QN => n1782);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3090, CK => CLK, Q => 
                           n_1685, QN => n1746);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3089, CK => CLK, Q => 
                           n_1686, QN => n1711);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3088, CK => CLK, Q => 
                           n_1687, QN => n1675);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3087, CK => CLK, Q => 
                           n_1688, QN => n1639);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3086, CK => CLK, Q => 
                           n_1689, QN => n1604);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3085, CK => CLK, Q => 
                           n_1690, QN => n1569);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3084, CK => CLK, Q => 
                           n_1691, QN => n1533);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3083, CK => CLK, Q => 
                           n_1692, QN => n1498);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3082, CK => CLK, Q => 
                           n_1693, QN => n1463);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3081, CK => CLK, Q => 
                           n_1694, QN => n1428);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3080, CK => CLK, Q => 
                           n_1695, QN => n1393);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3079, CK => CLK, Q => 
                           n_1696, QN => n1358);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3078, CK => CLK, Q => 
                           n_1697, QN => n1322);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3077, CK => CLK, Q => 
                           n_1698, QN => n1286);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3076, CK => CLK, Q => 
                           n_1699, QN => n1250);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3075, CK => CLK, Q => 
                           n_1700, QN => n1214);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3074, CK => CLK, Q => 
                           n_1701, QN => n1178);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3073, CK => CLK, Q => 
                           n_1702, QN => n1142);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3072, CK => CLK, Q => 
                           n_1703, QN => n1106);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3071, CK => CLK, Q => 
                           n_1704, QN => n1070);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3070, CK => CLK, Q => 
                           n_1705, QN => n2192);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3069, CK => CLK, Q => 
                           n_1706, QN => n2141);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3068, CK => CLK, Q => 
                           n_1707, QN => n2105);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3067, CK => CLK, Q => 
                           n_1708, QN => n2069);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3066, CK => CLK, Q => 
                           n_1709, QN => n2033);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3065, CK => CLK, Q => 
                           n_1710, QN => n1998);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3064, CK => CLK, Q => 
                           n_1711, QN => n1963);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3063, CK => CLK, Q => 
                           n_1712, QN => n1927);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3062, CK => CLK, Q => 
                           n_1713, QN => n1891);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3061, CK => CLK, Q => 
                           n_1714, QN => n1855);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3060, CK => CLK, Q => 
                           n_1715, QN => n1819);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3059, CK => CLK, Q => 
                           n_1716, QN => n1783);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3058, CK => CLK, Q => 
                           n_1717, QN => n1747);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3057, CK => CLK, Q => 
                           n_1718, QN => n1712);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3056, CK => CLK, Q => 
                           n_1719, QN => n1676);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3055, CK => CLK, Q => 
                           n_1720, QN => n1640);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3054, CK => CLK, Q => 
                           n_1721, QN => n1605);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3053, CK => CLK, Q => 
                           n_1722, QN => n1570);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3052, CK => CLK, Q => 
                           n_1723, QN => n1534);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3051, CK => CLK, Q => 
                           n_1724, QN => n1499);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3050, CK => CLK, Q => 
                           n_1725, QN => n1464);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3049, CK => CLK, Q => 
                           n_1726, QN => n1429);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3048, CK => CLK, Q => 
                           n_1727, QN => n1394);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3047, CK => CLK, Q => 
                           n_1728, QN => n1359);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => 
                           n_1729, QN => n1323);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => 
                           n_1730, QN => n1287);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => 
                           n_1731, QN => n1251);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => 
                           n_1732, QN => n1215);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => 
                           n_1733, QN => n1179);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => 
                           n_1734, QN => n1143);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => 
                           n_1735, QN => n1107);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => 
                           n_1736, QN => n1071);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => 
                           n3771, QN => n_1737);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => 
                           n3769, QN => n_1738);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => 
                           n3768, QN => n_1739);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => 
                           n3767, QN => n_1740);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => 
                           n3766, QN => n_1741);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => 
                           n3765, QN => n_1742);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => 
                           n3764, QN => n_1743);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => 
                           n3763, QN => n_1744);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => 
                           n3762, QN => n_1745);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => 
                           n3761, QN => n_1746);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => 
                           n3760, QN => n_1747);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => 
                           n3759, QN => n_1748);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => 
                           n3758, QN => n_1749);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => 
                           n3757, QN => n_1750);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => 
                           n3756, QN => n_1751);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => 
                           n3755, QN => n_1752);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => 
                           n3754, QN => n_1753);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => 
                           n3753, QN => n_1754);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => 
                           n3752, QN => n_1755);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => 
                           n3751, QN => n_1756);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => 
                           n3750, QN => n_1757);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => 
                           n3749, QN => n_1758);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => n3748
                           , QN => n_1759);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => n3747
                           , QN => n_1760);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => n3746
                           , QN => n_1761);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => n3745
                           , QN => n_1762);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => n3744
                           , QN => n_1763);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => n3743
                           , QN => n_1764);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => n3742
                           , QN => n_1765);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => n3741
                           , QN => n_1766);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => n3740
                           , QN => n_1767);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => n3739
                           , QN => n_1768);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => 
                           n3737, QN => n_1769);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => 
                           n3735, QN => n_1770);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => 
                           n3734, QN => n_1771);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => 
                           n3733, QN => n_1772);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => 
                           n3732, QN => n_1773);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => 
                           n3731, QN => n_1774);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => 
                           n3730, QN => n_1775);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => 
                           n3729, QN => n_1776);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => 
                           n3728, QN => n_1777);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => 
                           n3727, QN => n_1778);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => 
                           n3726, QN => n_1779);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => 
                           n3725, QN => n_1780);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => 
                           n3724, QN => n_1781);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => 
                           n3723, QN => n_1782);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => 
                           n3722, QN => n_1783);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => 
                           n3721, QN => n_1784);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => 
                           n3720, QN => n_1785);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => 
                           n3719, QN => n_1786);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => 
                           n3718, QN => n_1787);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => 
                           n3717, QN => n_1788);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => 
                           n3716, QN => n_1789);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => 
                           n3715, QN => n_1790);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => n3714
                           , QN => n_1791);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => n3713
                           , QN => n_1792);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n2982, CK => CLK, Q => n3712
                           , QN => n_1793);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n2981, CK => CLK, Q => n3711
                           , QN => n_1794);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n2980, CK => CLK, Q => n3710
                           , QN => n_1795);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n2979, CK => CLK, Q => n3709
                           , QN => n_1796);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n2978, CK => CLK, Q => n3708
                           , QN => n_1797);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n2977, CK => CLK, Q => n3707
                           , QN => n_1798);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n2976, CK => CLK, Q => n3706
                           , QN => n_1799);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n2975, CK => CLK, Q => n3705
                           , QN => n_1800);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n2974, CK => CLK, Q => 
                           n_1801, QN => n2185);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n2973, CK => CLK, Q => 
                           n_1802, QN => n2137);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n2972, CK => CLK, Q => 
                           n_1803, QN => n2101);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n2971, CK => CLK, Q => 
                           n_1804, QN => n2065);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n2970, CK => CLK, Q => 
                           n_1805, QN => n2029);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n2969, CK => CLK, Q => 
                           n_1806, QN => n1994);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n2968, CK => CLK, Q => 
                           n_1807, QN => n1959);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n2967, CK => CLK, Q => 
                           n_1808, QN => n1923);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n2966, CK => CLK, Q => 
                           n_1809, QN => n1887);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n2965, CK => CLK, Q => 
                           n_1810, QN => n1851);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n2964, CK => CLK, Q => 
                           n_1811, QN => n1815);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n2963, CK => CLK, Q => 
                           n_1812, QN => n1779);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n2962, CK => CLK, Q => 
                           n_1813, QN => n1743);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n2961, CK => CLK, Q => 
                           n_1814, QN => n1708);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n2960, CK => CLK, Q => 
                           n_1815, QN => n1672);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n2959, CK => CLK, Q => 
                           n_1816, QN => n1636);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n2958, CK => CLK, Q => 
                           n_1817, QN => n1601);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n2957, CK => CLK, Q => 
                           n_1818, QN => n1566);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n2956, CK => CLK, Q => 
                           n_1819, QN => n1530);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n2955, CK => CLK, Q => 
                           n_1820, QN => n1495);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n2954, CK => CLK, Q => 
                           n_1821, QN => n1460);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n2953, CK => CLK, Q => 
                           n_1822, QN => n1425);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n2952, CK => CLK, Q => 
                           n_1823, QN => n1390);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n2951, CK => CLK, Q => 
                           n_1824, QN => n1355);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n2950, CK => CLK, Q => 
                           n_1825, QN => n1319);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n2949, CK => CLK, Q => 
                           n_1826, QN => n1283);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n2948, CK => CLK, Q => 
                           n_1827, QN => n1247);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n2947, CK => CLK, Q => 
                           n_1828, QN => n1211);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n2946, CK => CLK, Q => 
                           n_1829, QN => n1175);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n2945, CK => CLK, Q => 
                           n_1830, QN => n1139);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n2944, CK => CLK, Q => 
                           n_1831, QN => n1103);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n2943, CK => CLK, Q => 
                           n_1832, QN => n1067);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n2942, CK => CLK, Q => 
                           n_1833, QN => n2187);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n2941, CK => CLK, Q => 
                           n_1834, QN => n2138);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n2940, CK => CLK, Q => 
                           n_1835, QN => n2102);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n2939, CK => CLK, Q => 
                           n_1836, QN => n2066);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n2938, CK => CLK, Q => 
                           n_1837, QN => n2030);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n2937, CK => CLK, Q => 
                           n_1838, QN => n1995);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n2936, CK => CLK, Q => 
                           n_1839, QN => n1960);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n2935, CK => CLK, Q => 
                           n_1840, QN => n1924);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n2934, CK => CLK, Q => 
                           n_1841, QN => n1888);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n2933, CK => CLK, Q => 
                           n_1842, QN => n1852);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n2932, CK => CLK, Q => 
                           n_1843, QN => n1816);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n2931, CK => CLK, Q => 
                           n_1844, QN => n1780);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n2930, CK => CLK, Q => 
                           n_1845, QN => n1744);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n2929, CK => CLK, Q => 
                           n_1846, QN => n1709);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n2928, CK => CLK, Q => 
                           n_1847, QN => n1673);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n2927, CK => CLK, Q => 
                           n_1848, QN => n1637);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n2926, CK => CLK, Q => 
                           n_1849, QN => n1602);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n2925, CK => CLK, Q => 
                           n_1850, QN => n1567);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n2924, CK => CLK, Q => 
                           n_1851, QN => n1531);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n2923, CK => CLK, Q => 
                           n_1852, QN => n1496);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n2922, CK => CLK, Q => 
                           n_1853, QN => n1461);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n2921, CK => CLK, Q => 
                           n_1854, QN => n1426);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n2920, CK => CLK, Q => 
                           n_1855, QN => n1391);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n2919, CK => CLK, Q => 
                           n_1856, QN => n1356);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n2918, CK => CLK, Q => 
                           n_1857, QN => n1320);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n2917, CK => CLK, Q => 
                           n_1858, QN => n1284);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n2916, CK => CLK, Q => 
                           n_1859, QN => n1248);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n2915, CK => CLK, Q => 
                           n_1860, QN => n1212);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n2914, CK => CLK, Q => 
                           n_1861, QN => n1176);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n2913, CK => CLK, Q => 
                           n_1862, QN => n1140);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n2912, CK => CLK, Q => 
                           n_1863, QN => n1104);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n2911, CK => CLK, Q => 
                           n_1864, QN => n1068);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n2910, CK => CLK, Q => 
                           n3635, QN => n_1865);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n2909, CK => CLK, Q => 
                           n3633, QN => n_1866);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n2908, CK => CLK, Q => 
                           n3632, QN => n_1867);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n2907, CK => CLK, Q => 
                           n3631, QN => n_1868);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n2906, CK => CLK, Q => 
                           n3630, QN => n_1869);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n2905, CK => CLK, Q => 
                           n3629, QN => n_1870);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n2904, CK => CLK, Q => 
                           n3628, QN => n_1871);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n2903, CK => CLK, Q => 
                           n3627, QN => n_1872);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n2902, CK => CLK, Q => 
                           n3626, QN => n_1873);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n2901, CK => CLK, Q => 
                           n3625, QN => n_1874);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n2900, CK => CLK, Q => 
                           n3624, QN => n_1875);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n2899, CK => CLK, Q => 
                           n3623, QN => n_1876);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n2898, CK => CLK, Q => 
                           n3622, QN => n_1877);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n2897, CK => CLK, Q => 
                           n3621, QN => n_1878);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n2896, CK => CLK, Q => 
                           n3620, QN => n_1879);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n2895, CK => CLK, Q => 
                           n3619, QN => n_1880);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n2894, CK => CLK, Q => 
                           n3618, QN => n_1881);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n2893, CK => CLK, Q => 
                           n3617, QN => n_1882);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n2892, CK => CLK, Q => 
                           n3616, QN => n_1883);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n2891, CK => CLK, Q => 
                           n3615, QN => n_1884);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n2890, CK => CLK, Q => 
                           n2526, QN => n_1885);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n2889, CK => CLK, Q => 
                           n2525, QN => n_1886);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n2888, CK => CLK, Q => n2524
                           , QN => n_1887);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n2887, CK => CLK, Q => n2523
                           , QN => n_1888);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n2886, CK => CLK, Q => n2522
                           , QN => n_1889);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n2885, CK => CLK, Q => n2521
                           , QN => n_1890);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n2884, CK => CLK, Q => n2520
                           , QN => n_1891);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n2883, CK => CLK, Q => n2519
                           , QN => n_1892);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n2882, CK => CLK, Q => n2518
                           , QN => n_1893);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n2881, CK => CLK, Q => n2517
                           , QN => n_1894);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n2880, CK => CLK, Q => n2516
                           , QN => n_1895);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n2879, CK => CLK, Q => n2515
                           , QN => n_1896);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n2878, CK => CLK, Q => 
                           n2513, QN => n_1897);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n2877, CK => CLK, Q => 
                           n2511, QN => n_1898);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n2876, CK => CLK, Q => 
                           n2510, QN => n_1899);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n2875, CK => CLK, Q => 
                           n2509, QN => n_1900);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n2874, CK => CLK, Q => 
                           n2508, QN => n_1901);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n2873, CK => CLK, Q => 
                           n2507, QN => n_1902);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n2872, CK => CLK, Q => 
                           n2506, QN => n_1903);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n2871, CK => CLK, Q => 
                           n2505, QN => n_1904);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n2870, CK => CLK, Q => 
                           n2504, QN => n_1905);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n2869, CK => CLK, Q => 
                           n2503, QN => n_1906);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n2868, CK => CLK, Q => 
                           n2502, QN => n_1907);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n2867, CK => CLK, Q => 
                           n2501, QN => n_1908);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n2866, CK => CLK, Q => 
                           n2500, QN => n_1909);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => 
                           n2499, QN => n_1910);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => 
                           n2498, QN => n_1911);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => 
                           n2497, QN => n_1912);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => 
                           n2496, QN => n_1913);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => 
                           n2495, QN => n_1914);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n2860, CK => CLK, Q => 
                           n2494, QN => n_1915);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n2859, CK => CLK, Q => 
                           n2493, QN => n_1916);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n2858, CK => CLK, Q => 
                           n2492, QN => n_1917);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n2857, CK => CLK, Q => 
                           n2491, QN => n_1918);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n2856, CK => CLK, Q => n2490
                           , QN => n_1919);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n2855, CK => CLK, Q => n2489
                           , QN => n_1920);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n2854, CK => CLK, Q => n2488
                           , QN => n_1921);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n2853, CK => CLK, Q => n2487
                           , QN => n_1922);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n2852, CK => CLK, Q => n2486
                           , QN => n_1923);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n2851, CK => CLK, Q => n2485
                           , QN => n_1924);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n2850, CK => CLK, Q => n2484
                           , QN => n_1925);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n2849, CK => CLK, Q => n2483
                           , QN => n_1926);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n2848, CK => CLK, Q => n2482
                           , QN => n_1927);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n2847, CK => CLK, Q => n2481
                           , QN => n_1928);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n2846, CK => CLK, Q => 
                           n2479, QN => n_1929);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n2845, CK => CLK, Q => 
                           n2477, QN => n_1930);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n2844, CK => CLK, Q => 
                           n2476, QN => n_1931);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n2843, CK => CLK, Q => 
                           n2475, QN => n_1932);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n2842, CK => CLK, Q => 
                           n2474, QN => n_1933);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n2841, CK => CLK, Q => 
                           n2473, QN => n_1934);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n2840, CK => CLK, Q => 
                           n2472, QN => n_1935);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => 
                           n2471, QN => n_1936);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n2838, CK => CLK, Q => 
                           n2470, QN => n_1937);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n2837, CK => CLK, Q => 
                           n2469, QN => n_1938);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n2836, CK => CLK, Q => 
                           n2468, QN => n_1939);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n2835, CK => CLK, Q => 
                           n2467, QN => n_1940);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n2834, CK => CLK, Q => 
                           n2466, QN => n_1941);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n2833, CK => CLK, Q => 
                           n2465, QN => n_1942);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n2832, CK => CLK, Q => 
                           n2464, QN => n_1943);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n2831, CK => CLK, Q => 
                           n2463, QN => n_1944);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n2830, CK => CLK, Q => 
                           n2462, QN => n_1945);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n2829, CK => CLK, Q => 
                           n2461, QN => n_1946);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n2828, CK => CLK, Q => 
                           n2460, QN => n_1947);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n2827, CK => CLK, Q => 
                           n2459, QN => n_1948);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n2826, CK => CLK, Q => 
                           n2458, QN => n_1949);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n2825, CK => CLK, Q => 
                           n2457, QN => n_1950);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n2824, CK => CLK, Q => n2456
                           , QN => n_1951);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n2823, CK => CLK, Q => n2455
                           , QN => n_1952);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n2822, CK => CLK, Q => n2454
                           , QN => n_1953);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n2821, CK => CLK, Q => n2453
                           , QN => n_1954);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n2820, CK => CLK, Q => n2452
                           , QN => n_1955);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n2819, CK => CLK, Q => n2451
                           , QN => n_1956);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n2818, CK => CLK, Q => n2450
                           , QN => n_1957);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n2817, CK => CLK, Q => n2449
                           , QN => n_1958);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n2816, CK => CLK, Q => n2448
                           , QN => n_1959);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n2815, CK => CLK, Q => n2447
                           , QN => n_1960);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n2814, CK => CLK, Q => 
                           n2441, QN => n_1961);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n2813, CK => CLK, Q => 
                           n2439, QN => n_1962);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n2812, CK => CLK, Q => 
                           n2438, QN => n_1963);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n2811, CK => CLK, Q => 
                           n2437, QN => n_1964);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n2810, CK => CLK, Q => 
                           n2436, QN => n_1965);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n2809, CK => CLK, Q => 
                           n2435, QN => n_1966);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n2808, CK => CLK, Q => 
                           n2434, QN => n_1967);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n2807, CK => CLK, Q => 
                           n2433, QN => n_1968);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n2806, CK => CLK, Q => 
                           n2432, QN => n_1969);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n2805, CK => CLK, Q => 
                           n2431, QN => n_1970);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n2804, CK => CLK, Q => 
                           n2430, QN => n_1971);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n2803, CK => CLK, Q => 
                           n2429, QN => n_1972);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n2802, CK => CLK, Q => 
                           n2428, QN => n_1973);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n2801, CK => CLK, Q => 
                           n2427, QN => n_1974);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n2800, CK => CLK, Q => 
                           n2426, QN => n_1975);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n2799, CK => CLK, Q => 
                           n2425, QN => n_1976);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n2798, CK => CLK, Q => 
                           n2424, QN => n_1977);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n2797, CK => CLK, Q => 
                           n2423, QN => n_1978);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n2796, CK => CLK, Q => 
                           n2422, QN => n_1979);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n2795, CK => CLK, Q => 
                           n2421, QN => n_1980);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n2794, CK => CLK, Q => 
                           n2420, QN => n_1981);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n2793, CK => CLK, Q => 
                           n2419, QN => n_1982);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n2792, CK => CLK, Q => n2418
                           , QN => n_1983);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n2791, CK => CLK, Q => n2417
                           , QN => n_1984);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n2790, CK => CLK, Q => n2416
                           , QN => n_1985);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n2789, CK => CLK, Q => n2415
                           , QN => n_1986);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n2788, CK => CLK, Q => n2414
                           , QN => n_1987);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n2787, CK => CLK, Q => n2413
                           , QN => n_1988);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n2786, CK => CLK, Q => n2412
                           , QN => n_1989);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n2785, CK => CLK, Q => n2411
                           , QN => n_1990);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n2784, CK => CLK, Q => n2410
                           , QN => n_1991);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n2783, CK => CLK, Q => n2409
                           , QN => n_1992);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n2782, CK => CLK, Q => 
                           n_1993, QN => n2180);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n2781, CK => CLK, Q => 
                           n_1994, QN => n2134);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n2780, CK => CLK, Q => 
                           n_1995, QN => n2098);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n2779, CK => CLK, Q => 
                           n_1996, QN => n2062);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n2778, CK => CLK, Q => 
                           n_1997, QN => n2026);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n2777, CK => CLK, Q => 
                           n_1998, QN => n1991);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n2776, CK => CLK, Q => 
                           n_1999, QN => n1956);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n2775, CK => CLK, Q => 
                           n_2000, QN => n1920);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n2774, CK => CLK, Q => 
                           n_2001, QN => n1884);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n2773, CK => CLK, Q => 
                           n_2002, QN => n1848);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n2772, CK => CLK, Q => 
                           n_2003, QN => n1812);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n2771, CK => CLK, Q => 
                           n_2004, QN => n1776);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n2770, CK => CLK, Q => 
                           n_2005, QN => n1740);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n2769, CK => CLK, Q => 
                           n_2006, QN => n1705);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n2768, CK => CLK, Q => 
                           n_2007, QN => n1669);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n2767, CK => CLK, Q => 
                           n_2008, QN => n1633);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n2766, CK => CLK, Q => 
                           n_2009, QN => n1598);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n2765, CK => CLK, Q => 
                           n_2010, QN => n1563);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n2764, CK => CLK, Q => 
                           n_2011, QN => n1527);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n2763, CK => CLK, Q => 
                           n_2012, QN => n1492);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n2762, CK => CLK, Q => 
                           n_2013, QN => n1457);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n2761, CK => CLK, Q => 
                           n_2014, QN => n1422);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n2760, CK => CLK, Q => 
                           n_2015, QN => n1387);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n2759, CK => CLK, Q => 
                           n_2016, QN => n1352);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n2758, CK => CLK, Q => 
                           n_2017, QN => n1316);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n2757, CK => CLK, Q => 
                           n_2018, QN => n1280);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n2756, CK => CLK, Q => 
                           n_2019, QN => n1244);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n2755, CK => CLK, Q => 
                           n_2020, QN => n1208);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n2754, CK => CLK, Q => 
                           n_2021, QN => n1172);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n2753, CK => CLK, Q => 
                           n_2022, QN => n1136);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n2752, CK => CLK, Q => 
                           n_2023, QN => n1100);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n2751, CK => CLK, Q => 
                           n_2024, QN => n1062);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n2750, CK => CLK, Q => 
                           n_2025, QN => n2182);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n2749, CK => CLK, Q => 
                           n_2026, QN => n2135);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n2748, CK => CLK, Q => 
                           n_2027, QN => n2099);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n2747, CK => CLK, Q => 
                           n_2028, QN => n2063);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n2746, CK => CLK, Q => 
                           n_2029, QN => n2027);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n2745, CK => CLK, Q => 
                           n_2030, QN => n1992);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n2744, CK => CLK, Q => 
                           n_2031, QN => n1957);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n2743, CK => CLK, Q => 
                           n_2032, QN => n1921);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n2742, CK => CLK, Q => 
                           n_2033, QN => n1885);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n2741, CK => CLK, Q => 
                           n_2034, QN => n1849);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n2740, CK => CLK, Q => 
                           n_2035, QN => n1813);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n2739, CK => CLK, Q => 
                           n_2036, QN => n1777);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n2738, CK => CLK, Q => 
                           n_2037, QN => n1741);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n2737, CK => CLK, Q => 
                           n_2038, QN => n1706);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n2736, CK => CLK, Q => 
                           n_2039, QN => n1670);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n2735, CK => CLK, Q => 
                           n_2040, QN => n1634);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n2734, CK => CLK, Q => 
                           n_2041, QN => n1599);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n2733, CK => CLK, Q => 
                           n_2042, QN => n1564);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n2732, CK => CLK, Q => 
                           n_2043, QN => n1528);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n2731, CK => CLK, Q => 
                           n_2044, QN => n1493);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n2730, CK => CLK, Q => 
                           n_2045, QN => n1458);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n2729, CK => CLK, Q => 
                           n_2046, QN => n1423);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n2728, CK => CLK, Q => 
                           n_2047, QN => n1388);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n2727, CK => CLK, Q => 
                           n_2048, QN => n1353);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n2726, CK => CLK, Q => 
                           n_2049, QN => n1317);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n2725, CK => CLK, Q => 
                           n_2050, QN => n1281);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n2724, CK => CLK, Q => 
                           n_2051, QN => n1245);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n2723, CK => CLK, Q => 
                           n_2052, QN => n1209);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n2722, CK => CLK, Q => 
                           n_2053, QN => n1173);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n2721, CK => CLK, Q => 
                           n_2054, QN => n1137);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n2720, CK => CLK, Q => 
                           n_2055, QN => n1101);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n2719, CK => CLK, Q => 
                           n_2056, QN => n1063);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n2718, CK => CLK, Q => 
                           n2339, QN => n_2057);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n2717, CK => CLK, Q => 
                           n2337, QN => n_2058);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n2716, CK => CLK, Q => 
                           n2336, QN => n_2059);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n2715, CK => CLK, Q => 
                           n2335, QN => n_2060);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n2714, CK => CLK, Q => 
                           n2334, QN => n_2061);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n2713, CK => CLK, Q => 
                           n2333, QN => n_2062);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n2712, CK => CLK, Q => 
                           n2332, QN => n_2063);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n2711, CK => CLK, Q => 
                           n2331, QN => n_2064);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n2710, CK => CLK, Q => 
                           n2330, QN => n_2065);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n2709, CK => CLK, Q => 
                           n2329, QN => n_2066);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n2708, CK => CLK, Q => 
                           n2328, QN => n_2067);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n2707, CK => CLK, Q => 
                           n2327, QN => n_2068);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n2706, CK => CLK, Q => 
                           n2326, QN => n_2069);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n2705, CK => CLK, Q => 
                           n2325, QN => n_2070);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n2704, CK => CLK, Q => 
                           n2324, QN => n_2071);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n2703, CK => CLK, Q => 
                           n2323, QN => n_2072);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n2702, CK => CLK, Q => 
                           n2322, QN => n_2073);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n2701, CK => CLK, Q => 
                           n2321, QN => n_2074);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n2700, CK => CLK, Q => 
                           n2320, QN => n_2075);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n2699, CK => CLK, Q => 
                           n2319, QN => n_2076);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n2698, CK => CLK, Q => 
                           n2318, QN => n_2077);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n2697, CK => CLK, Q => 
                           n2317, QN => n_2078);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n2696, CK => CLK, Q => n2316
                           , QN => n_2079);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n2695, CK => CLK, Q => n2315
                           , QN => n_2080);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n2694, CK => CLK, Q => n2314
                           , QN => n_2081);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n2693, CK => CLK, Q => n2313
                           , QN => n_2082);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n2692, CK => CLK, Q => n2312
                           , QN => n_2083);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n2691, CK => CLK, Q => n2311
                           , QN => n_2084);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n2690, CK => CLK, Q => n2310
                           , QN => n_2085);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n2689, CK => CLK, Q => n2309
                           , QN => n_2086);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n2688, CK => CLK, Q => n2308
                           , QN => n_2087);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n2687, CK => CLK, Q => n2307
                           , QN => n_2088);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n2686, CK => CLK, Q => 
                           n2305, QN => n_2089);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n2685, CK => CLK, Q => 
                           n2303, QN => n_2090);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n2684, CK => CLK, Q => 
                           n2302, QN => n_2091);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n2683, CK => CLK, Q => 
                           n2301, QN => n_2092);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n2682, CK => CLK, Q => 
                           n2300, QN => n_2093);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n2681, CK => CLK, Q => 
                           n2299, QN => n_2094);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n2680, CK => CLK, Q => 
                           n2298, QN => n_2095);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n2679, CK => CLK, Q => 
                           n2297, QN => n_2096);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n2678, CK => CLK, Q => 
                           n2296, QN => n_2097);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n2677, CK => CLK, Q => 
                           n2295, QN => n_2098);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n2676, CK => CLK, Q => 
                           n2294, QN => n_2099);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n2675, CK => CLK, Q => 
                           n2293, QN => n_2100);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n2674, CK => CLK, Q => 
                           n2292, QN => n_2101);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n2673, CK => CLK, Q => 
                           n2291, QN => n_2102);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n2672, CK => CLK, Q => 
                           n2290, QN => n_2103);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n2671, CK => CLK, Q => 
                           n2289, QN => n_2104);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n2670, CK => CLK, Q => 
                           n2288, QN => n_2105);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n2669, CK => CLK, Q => 
                           n2287, QN => n_2106);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n2668, CK => CLK, Q => 
                           n2286, QN => n_2107);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n2667, CK => CLK, Q => 
                           n2285, QN => n_2108);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n2666, CK => CLK, Q => 
                           n2284, QN => n_2109);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n2665, CK => CLK, Q => 
                           n2283, QN => n_2110);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n2664, CK => CLK, Q => n2282
                           , QN => n_2111);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n2663, CK => CLK, Q => n2281
                           , QN => n_2112);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n2662, CK => CLK, Q => n2280
                           , QN => n_2113);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n2661, CK => CLK, Q => n2279
                           , QN => n_2114);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n2660, CK => CLK, Q => n2278
                           , QN => n_2115);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n2659, CK => CLK, Q => n2277
                           , QN => n_2116);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n2658, CK => CLK, Q => n2276
                           , QN => n_2117);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n2657, CK => CLK, Q => n2275
                           , QN => n_2118);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n2656, CK => CLK, Q => n2274
                           , QN => n_2119);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n2655, CK => CLK, Q => n2273
                           , QN => n_2120);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n2654, CK => CLK, Q => 
                           n_2121, QN => n2175);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n2653, CK => CLK, Q => 
                           n_2122, QN => n2131);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n2652, CK => CLK, Q => 
                           n_2123, QN => n2095);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n2651, CK => CLK, Q => 
                           n_2124, QN => n2059);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n2650, CK => CLK, Q => 
                           n_2125, QN => n2023);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n2649, CK => CLK, Q => 
                           n_2126, QN => n1988);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n2648, CK => CLK, Q => 
                           n_2127, QN => n1953);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n2647, CK => CLK, Q => 
                           n_2128, QN => n1917);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n2646, CK => CLK, Q => 
                           n_2129, QN => n1881);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n2645, CK => CLK, Q => 
                           n_2130, QN => n1845);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n2644, CK => CLK, Q => 
                           n_2131, QN => n1809);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n2643, CK => CLK, Q => 
                           n_2132, QN => n1773);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n2642, CK => CLK, Q => 
                           n_2133, QN => n1737);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n2641, CK => CLK, Q => 
                           n_2134, QN => n1702);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n2640, CK => CLK, Q => 
                           n_2135, QN => n1666);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n2639, CK => CLK, Q => 
                           n_2136, QN => n1630);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n2638, CK => CLK, Q => 
                           n_2137, QN => n1595);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n2637, CK => CLK, Q => 
                           n_2138, QN => n1560);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n2636, CK => CLK, Q => 
                           n_2139, QN => n1524);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n2635, CK => CLK, Q => 
                           n_2140, QN => n1489);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n2634, CK => CLK, Q => 
                           n_2141, QN => n1454);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n2633, CK => CLK, Q => 
                           n_2142, QN => n1419);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n2632, CK => CLK, Q => 
                           n_2143, QN => n1384);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n2631, CK => CLK, Q => 
                           n_2144, QN => n1349);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n2630, CK => CLK, Q => 
                           n_2145, QN => n1313);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n2629, CK => CLK, Q => 
                           n_2146, QN => n1277);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n2628, CK => CLK, Q => 
                           n_2147, QN => n1241);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n2627, CK => CLK, Q => 
                           n_2148, QN => n1205);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n2626, CK => CLK, Q => 
                           n_2149, QN => n1169);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n2625, CK => CLK, Q => 
                           n_2150, QN => n1133);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n2624, CK => CLK, Q => 
                           n_2151, QN => n1097);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n2623, CK => CLK, Q => 
                           n_2152, QN => n1059);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n2622, CK => CLK, Q => 
                           n_2153, QN => n2177);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n2621, CK => CLK, Q => 
                           n_2154, QN => n2132);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n2620, CK => CLK, Q => 
                           n_2155, QN => n2096);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n2619, CK => CLK, Q => 
                           n_2156, QN => n2060);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n2618, CK => CLK, Q => 
                           n_2157, QN => n2024);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n2617, CK => CLK, Q => 
                           n_2158, QN => n1989);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n2616, CK => CLK, Q => 
                           n_2159, QN => n1954);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n2615, CK => CLK, Q => 
                           n_2160, QN => n1918);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n2614, CK => CLK, Q => 
                           n_2161, QN => n1882);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n2613, CK => CLK, Q => 
                           n_2162, QN => n1846);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n2612, CK => CLK, Q => 
                           n_2163, QN => n1810);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n2611, CK => CLK, Q => 
                           n_2164, QN => n1774);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n2610, CK => CLK, Q => 
                           n_2165, QN => n1738);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n2609, CK => CLK, Q => 
                           n_2166, QN => n1703);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n2608, CK => CLK, Q => 
                           n_2167, QN => n1667);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n2607, CK => CLK, Q => 
                           n_2168, QN => n1631);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n2606, CK => CLK, Q => 
                           n_2169, QN => n1596);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n2605, CK => CLK, Q => 
                           n_2170, QN => n1561);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n2604, CK => CLK, Q => 
                           n_2171, QN => n1525);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n2603, CK => CLK, Q => 
                           n_2172, QN => n1490);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n2602, CK => CLK, Q => 
                           n_2173, QN => n1455);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n2601, CK => CLK, Q => 
                           n_2174, QN => n1420);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n2600, CK => CLK, Q => 
                           n_2175, QN => n1385);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n2599, CK => CLK, Q => 
                           n_2176, QN => n1350);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n2598, CK => CLK, Q => 
                           n_2177, QN => n1314);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n2597, CK => CLK, Q => 
                           n_2178, QN => n1278);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n2596, CK => CLK, Q => 
                           n_2179, QN => n1242);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n2595, CK => CLK, Q => 
                           n_2180, QN => n1206);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n2594, CK => CLK, Q => 
                           n_2181, QN => n1170);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n2593, CK => CLK, Q => 
                           n_2182, QN => n1134);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n2592, CK => CLK, Q => 
                           n_2183, QN => n1098);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n2591, CK => CLK, Q => 
                           n_2184, QN => n1060);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2582, CK => CLK, Q => OUT1(23), QN
                           => n1900);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2581, CK => CLK, Q => OUT1(22), QN
                           => n1864);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2580, CK => CLK, Q => OUT1(21), QN
                           => n1828);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2579, CK => CLK, Q => OUT1(20), QN
                           => n1792);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2578, CK => CLK, Q => OUT1(19), QN
                           => n1756);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2577, CK => CLK, Q => OUT1(18), QN
                           => n17);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2576, CK => CLK, Q => OUT1(17), QN
                           => n1685);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2575, CK => CLK, Q => OUT1(16), QN
                           => n1649);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2574, CK => CLK, Q => OUT1(15), QN
                           => n22);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2573, CK => CLK, Q => OUT1(14), QN
                           => n21);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2572, CK => CLK, Q => OUT1(13), QN
                           => n1543);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2571, CK => CLK, Q => OUT1(12), QN
                           => n25);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2570, CK => CLK, Q => OUT1(11), QN
                           => n24);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => OUT1(5), QN 
                           => n1260);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => OUT1(4), QN 
                           => n1224);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => OUT1(3), QN 
                           => n1188);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => OUT1(2), QN 
                           => n1152);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => OUT1(1), QN 
                           => n1116);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => OUT1(0), QN 
                           => n1080);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => OUT2(23), QN
                           => n864);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => OUT2(22), QN
                           => n844);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => OUT2(21), QN
                           => n13);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => OUT2(20), QN
                           => n805);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => OUT2(19), QN
                           => n785);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => OUT2(18), QN
                           => n11);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => OUT2(17), QN
                           => n10);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => OUT2(16), QN
                           => n727);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => OUT2(15), QN
                           => n707);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => OUT2(14), QN
                           => n18);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => OUT2(13), QN
                           => n668);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => OUT2(12), QN
                           => n648);
   U3 : AND2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1);
   U4 : AND2_X1 port map( A1 => ADD_RD2(1), A2 => n391, ZN => n2);
   U5 : AND2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n3);
   U6 : AND2_X1 port map( A1 => ADD_RD1(1), A2 => n1043, ZN => n4);
   U7 : AND2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), ZN => n15);
   U8 : AND2_X1 port map( A1 => ADD_WR(4), A2 => WR, ZN => n16);
   U9 : CLKBUF_X3 port map( A => n2203, Z => n291);
   U10 : CLKBUF_X3 port map( A => n1039, Z => n189);
   U11 : BUF_X1 port map( A => n2167, Z => n229);
   U12 : BUF_X1 port map( A => n1012, Z => n127);
   U13 : BUF_X2 port map( A => n1019, Z => n139);
   U14 : BUF_X2 port map( A => n1003, Z => n91);
   U15 : BUF_X2 port map( A => n1023, Z => n154);
   U16 : BUF_X2 port map( A => n1029, Z => n178);
   U17 : BUF_X2 port map( A => n1026, Z => n166);
   U18 : BUF_X2 port map( A => n1007, Z => n106);
   U19 : BUF_X2 port map( A => n1013, Z => n130);
   U20 : BUF_X2 port map( A => n1010, Z => n118);
   U21 : BUF_X2 port map( A => n1004, Z => n94);
   U22 : BUF_X1 port map( A => n2193, Z => n279);
   U23 : BUF_X1 port map( A => n2193, Z => n280);
   U24 : BUF_X1 port map( A => n2188, Z => n267);
   U25 : BUF_X1 port map( A => n2188, Z => n268);
   U26 : BUF_X1 port map( A => n2159, Z => n208);
   U27 : BUF_X1 port map( A => n2169, Z => n232);
   U28 : BUF_X1 port map( A => n2164, Z => n220);
   U29 : BUF_X1 port map( A => n2154, Z => n196);
   U30 : BUF_X1 port map( A => n2178, Z => n243);
   U31 : BUF_X1 port map( A => n2178, Z => n244);
   U32 : BUF_X1 port map( A => n2181, Z => n252);
   U33 : BUF_X1 port map( A => n2181, Z => n253);
   U34 : BUF_X1 port map( A => n2186, Z => n264);
   U35 : BUF_X1 port map( A => n2186, Z => n265);
   U36 : BUF_X1 port map( A => n2191, Z => n276);
   U37 : BUF_X1 port map( A => n2191, Z => n277);
   U38 : BUF_X1 port map( A => n2157, Z => n205);
   U39 : BUF_X1 port map( A => n2162, Z => n217);
   U40 : BUF_X1 port map( A => n2176, Z => n240);
   U41 : BUF_X1 port map( A => n2176, Z => n241);
   U42 : BUF_X1 port map( A => n2152, Z => n193);
   U43 : BUF_X1 port map( A => n1022, Z => n151);
   U44 : BUF_X1 port map( A => n1025, Z => n163);
   U45 : BUF_X1 port map( A => n1028, Z => n175);
   U46 : BUF_X1 port map( A => n1006, Z => n103);
   U47 : BUF_X1 port map( A => n1009, Z => n115);
   U48 : BUF_X1 port map( A => n1039, Z => n191);
   U49 : BUF_X1 port map( A => n2203, Z => n293);
   U50 : BUF_X2 port map( A => n2270, Z => n297);
   U51 : BUF_X2 port map( A => n2270, Z => n298);
   U52 : BUF_X2 port map( A => n2372, Z => n306);
   U53 : BUF_X2 port map( A => n2372, Z => n307);
   U54 : BUF_X2 port map( A => n2406, Z => n309);
   U55 : BUF_X2 port map( A => n2406, Z => n310);
   U56 : BUF_X2 port map( A => n3804, Z => n336);
   U57 : BUF_X2 port map( A => n3804, Z => n337);
   U58 : BUF_X2 port map( A => n3839, Z => n339);
   U59 : BUF_X2 port map( A => n3839, Z => n340);
   U60 : BUF_X2 port map( A => n2236, Z => n294);
   U61 : BUF_X2 port map( A => n2236, Z => n295);
   U62 : BUF_X2 port map( A => n3668, Z => n324);
   U63 : BUF_X2 port map( A => n3668, Z => n325);
   U64 : BUF_X2 port map( A => n3702, Z => n327);
   U65 : BUF_X2 port map( A => n3702, Z => n328);
   U66 : BUF_X2 port map( A => n2304, Z => n300);
   U67 : BUF_X2 port map( A => n2304, Z => n301);
   U68 : BUF_X2 port map( A => n2338, Z => n303);
   U69 : BUF_X2 port map( A => n2338, Z => n304);
   U70 : BUF_X2 port map( A => n2440, Z => n312);
   U71 : BUF_X2 port map( A => n2440, Z => n313);
   U72 : BUF_X2 port map( A => n2478, Z => n315);
   U73 : BUF_X2 port map( A => n2478, Z => n316);
   U74 : BUF_X2 port map( A => n2512, Z => n318);
   U75 : BUF_X2 port map( A => n2512, Z => n319);
   U76 : BUF_X2 port map( A => n3736, Z => n330);
   U77 : BUF_X2 port map( A => n3736, Z => n331);
   U78 : BUF_X2 port map( A => n3634, Z => n321);
   U79 : BUF_X2 port map( A => n3634, Z => n322);
   U80 : BUF_X2 port map( A => n3770, Z => n333);
   U81 : BUF_X2 port map( A => n3770, Z => n334);
   U82 : BUF_X1 port map( A => n27, Z => n288);
   U83 : BUF_X1 port map( A => n28, Z => n186);
   U84 : BUF_X1 port map( A => n28, Z => n187);
   U85 : BUF_X1 port map( A => n27, Z => n289);
   U86 : BUF_X2 port map( A => n2167, Z => n228);
   U87 : BUF_X1 port map( A => n29, Z => n156);
   U88 : BUF_X1 port map( A => n29, Z => n157);
   U89 : BUF_X1 port map( A => n30, Z => n258);
   U90 : BUF_X1 port map( A => n30, Z => n259);
   U91 : BUF_X2 port map( A => n1012, Z => n126);
   U92 : BUF_X1 port map( A => n2270, Z => n299);
   U93 : BUF_X1 port map( A => n2372, Z => n308);
   U94 : BUF_X1 port map( A => n2406, Z => n311);
   U95 : BUF_X1 port map( A => n3804, Z => n338);
   U96 : BUF_X1 port map( A => n3839, Z => n341);
   U97 : BUF_X1 port map( A => n2236, Z => n296);
   U98 : BUF_X1 port map( A => n3668, Z => n326);
   U99 : BUF_X1 port map( A => n3702, Z => n329);
   U100 : BUF_X1 port map( A => n2304, Z => n302);
   U101 : BUF_X1 port map( A => n2338, Z => n305);
   U102 : BUF_X1 port map( A => n2440, Z => n314);
   U103 : BUF_X1 port map( A => n2478, Z => n317);
   U104 : BUF_X1 port map( A => n2512, Z => n320);
   U105 : BUF_X1 port map( A => n3736, Z => n332);
   U106 : BUF_X1 port map( A => n3634, Z => n323);
   U107 : BUF_X1 port map( A => n3770, Z => n335);
   U108 : BUF_X1 port map( A => n28, Z => n188);
   U109 : BUF_X1 port map( A => n27, Z => n290);
   U110 : BUF_X1 port map( A => n2167, Z => n230);
   U111 : BUF_X1 port map( A => n29, Z => n158);
   U112 : BUF_X1 port map( A => n30, Z => n260);
   U113 : BUF_X1 port map( A => n1012, Z => n128);
   U114 : BUF_X2 port map( A => n3941, Z => n348);
   U115 : BUF_X2 port map( A => n3941, Z => n349);
   U116 : BUF_X2 port map( A => n3975, Z => n351);
   U117 : BUF_X2 port map( A => n3975, Z => n352);
   U118 : BUF_X2 port map( A => n4077, Z => n360);
   U119 : BUF_X2 port map( A => n4077, Z => n361);
   U120 : BUF_X2 port map( A => n4112, Z => n363);
   U121 : BUF_X2 port map( A => n4112, Z => n364);
   U122 : BUF_X2 port map( A => n4458, Z => n387);
   U123 : BUF_X2 port map( A => n4458, Z => n388);
   U124 : BUF_X2 port map( A => n4219, Z => n372);
   U125 : BUF_X2 port map( A => n4219, Z => n373);
   U126 : BUF_X2 port map( A => n4254, Z => n375);
   U127 : BUF_X2 port map( A => n4254, Z => n376);
   U128 : BUF_X2 port map( A => n4391, Z => n384);
   U129 : BUF_X2 port map( A => n4391, Z => n385);
   U130 : BUF_X2 port map( A => n3873, Z => n342);
   U131 : BUF_X2 port map( A => n3873, Z => n343);
   U132 : BUF_X2 port map( A => n3907, Z => n345);
   U133 : BUF_X2 port map( A => n3907, Z => n346);
   U134 : BUF_X2 port map( A => n4009, Z => n354);
   U135 : BUF_X2 port map( A => n4009, Z => n355);
   U136 : BUF_X2 port map( A => n4043, Z => n357);
   U137 : BUF_X2 port map( A => n4043, Z => n358);
   U138 : BUF_X2 port map( A => n4184, Z => n369);
   U139 : BUF_X2 port map( A => n4184, Z => n370);
   U140 : BUF_X2 port map( A => n4149, Z => n366);
   U141 : BUF_X2 port map( A => n4149, Z => n367);
   U142 : BUF_X2 port map( A => n4289, Z => n378);
   U143 : BUF_X2 port map( A => n4289, Z => n379);
   U144 : BUF_X2 port map( A => n4355, Z => n381);
   U145 : BUF_X2 port map( A => n4355, Z => n382);
   U146 : BUF_X2 port map( A => n2159, Z => n207);
   U147 : BUF_X2 port map( A => n2164, Z => n219);
   U148 : BUF_X2 port map( A => n2169, Z => n231);
   U149 : BUF_X2 port map( A => n2154, Z => n195);
   U150 : BUF_X2 port map( A => n2183, Z => n255);
   U151 : BUF_X2 port map( A => n2183, Z => n256);
   U152 : BUF_X2 port map( A => n2157, Z => n204);
   U153 : BUF_X2 port map( A => n2162, Z => n216);
   U154 : BUF_X2 port map( A => n2152, Z => n192);
   U155 : BUF_X1 port map( A => n47, Z => n210);
   U156 : BUF_X1 port map( A => n48, Z => n222);
   U157 : BUF_X1 port map( A => n50, Z => n234);
   U158 : BUF_X1 port map( A => n54, Z => n198);
   U159 : BUF_X1 port map( A => n49, Z => n168);
   U160 : BUF_X1 port map( A => n51, Z => n180);
   U161 : BUF_X1 port map( A => n52, Z => n108);
   U162 : BUF_X1 port map( A => n53, Z => n120);
   U163 : BUF_X1 port map( A => n55, Z => n132);
   U164 : BUF_X1 port map( A => n41, Z => n144);
   U165 : BUF_X1 port map( A => n56, Z => n96);
   U166 : BUF_X1 port map( A => n59, Z => n270);
   U167 : BUF_X1 port map( A => n60, Z => n282);
   U168 : BUF_X1 port map( A => n42, Z => n246);
   U169 : BUF_X1 port map( A => n49, Z => n169);
   U170 : BUF_X1 port map( A => n51, Z => n181);
   U171 : BUF_X1 port map( A => n52, Z => n109);
   U172 : BUF_X1 port map( A => n53, Z => n121);
   U173 : BUF_X1 port map( A => n55, Z => n133);
   U174 : BUF_X1 port map( A => n41, Z => n145);
   U175 : BUF_X1 port map( A => n59, Z => n271);
   U176 : BUF_X1 port map( A => n56, Z => n97);
   U177 : BUF_X1 port map( A => n60, Z => n283);
   U178 : BUF_X1 port map( A => n47, Z => n211);
   U179 : BUF_X1 port map( A => n48, Z => n223);
   U180 : BUF_X1 port map( A => n50, Z => n235);
   U181 : BUF_X1 port map( A => n42, Z => n247);
   U182 : BUF_X1 port map( A => n54, Z => n199);
   U183 : BUF_X2 port map( A => n1025, Z => n162);
   U184 : BUF_X2 port map( A => n1028, Z => n174);
   U185 : BUF_X2 port map( A => n1006, Z => n102);
   U186 : BUF_X2 port map( A => n1009, Z => n114);
   U187 : BUF_X2 port map( A => n1003, Z => n90);
   U188 : BUF_X2 port map( A => n1022, Z => n150);
   U189 : BUF_X2 port map( A => n1019, Z => n138);
   U190 : BUF_X2 port map( A => n1026, Z => n165);
   U191 : BUF_X2 port map( A => n1029, Z => n177);
   U192 : BUF_X2 port map( A => n1007, Z => n105);
   U193 : BUF_X2 port map( A => n1010, Z => n117);
   U194 : BUF_X2 port map( A => n1013, Z => n129);
   U195 : BUF_X2 port map( A => n1004, Z => n93);
   U196 : BUF_X2 port map( A => n1023, Z => n153);
   U197 : BUF_X2 port map( A => n1020, Z => n141);
   U198 : BUF_X1 port map( A => n1020, Z => n142);
   U199 : BUF_X1 port map( A => n63, Z => n213);
   U200 : BUF_X1 port map( A => n61, Z => n225);
   U201 : BUF_X1 port map( A => n64, Z => n237);
   U202 : BUF_X1 port map( A => n45, Z => n201);
   U203 : BUF_X1 port map( A => n43, Z => n171);
   U204 : BUF_X1 port map( A => n44, Z => n183);
   U205 : BUF_X1 port map( A => n39, Z => n159);
   U206 : BUF_X1 port map( A => n65, Z => n111);
   U207 : BUF_X1 port map( A => n62, Z => n123);
   U208 : BUF_X1 port map( A => n66, Z => n135);
   U209 : BUF_X1 port map( A => n37, Z => n147);
   U210 : BUF_X1 port map( A => n46, Z => n99);
   U211 : BUF_X1 port map( A => n57, Z => n273);
   U212 : BUF_X1 port map( A => n58, Z => n285);
   U213 : BUF_X1 port map( A => n38, Z => n249);
   U214 : BUF_X1 port map( A => n43, Z => n172);
   U215 : BUF_X1 port map( A => n44, Z => n184);
   U216 : BUF_X1 port map( A => n39, Z => n160);
   U217 : BUF_X1 port map( A => n65, Z => n112);
   U218 : BUF_X1 port map( A => n62, Z => n124);
   U219 : BUF_X1 port map( A => n66, Z => n136);
   U220 : BUF_X1 port map( A => n37, Z => n148);
   U221 : BUF_X1 port map( A => n46, Z => n100);
   U222 : BUF_X1 port map( A => n57, Z => n274);
   U223 : BUF_X1 port map( A => n40, Z => n261);
   U224 : BUF_X1 port map( A => n40, Z => n262);
   U225 : BUF_X1 port map( A => n58, Z => n286);
   U226 : BUF_X1 port map( A => n63, Z => n214);
   U227 : BUF_X1 port map( A => n61, Z => n226);
   U228 : BUF_X1 port map( A => n38, Z => n250);
   U229 : BUF_X1 port map( A => n64, Z => n238);
   U230 : BUF_X1 port map( A => n45, Z => n202);
   U231 : BUF_X1 port map( A => n3941, Z => n350);
   U232 : BUF_X1 port map( A => n3975, Z => n353);
   U233 : BUF_X1 port map( A => n4077, Z => n362);
   U234 : BUF_X1 port map( A => n4112, Z => n365);
   U235 : BUF_X1 port map( A => n4458, Z => n389);
   U236 : BUF_X1 port map( A => n4219, Z => n374);
   U237 : BUF_X1 port map( A => n4254, Z => n377);
   U238 : BUF_X1 port map( A => n4391, Z => n386);
   U239 : BUF_X1 port map( A => n3873, Z => n344);
   U240 : BUF_X1 port map( A => n3907, Z => n347);
   U241 : BUF_X1 port map( A => n4009, Z => n356);
   U242 : BUF_X1 port map( A => n4043, Z => n359);
   U243 : BUF_X1 port map( A => n4184, Z => n371);
   U244 : BUF_X1 port map( A => n4149, Z => n368);
   U245 : BUF_X1 port map( A => n4289, Z => n380);
   U246 : BUF_X1 port map( A => n4355, Z => n383);
   U247 : BUF_X1 port map( A => n2188, Z => n269);
   U248 : BUF_X1 port map( A => n2193, Z => n281);
   U249 : BUF_X1 port map( A => n2159, Z => n209);
   U250 : BUF_X1 port map( A => n2164, Z => n221);
   U251 : BUF_X1 port map( A => n2169, Z => n233);
   U252 : BUF_X1 port map( A => n2154, Z => n197);
   U253 : BUF_X1 port map( A => n2183, Z => n257);
   U254 : BUF_X1 port map( A => n2178, Z => n245);
   U255 : BUF_X1 port map( A => n2186, Z => n266);
   U256 : BUF_X1 port map( A => n2191, Z => n278);
   U257 : BUF_X1 port map( A => n2157, Z => n206);
   U258 : BUF_X1 port map( A => n2162, Z => n218);
   U259 : BUF_X1 port map( A => n2152, Z => n194);
   U260 : BUF_X1 port map( A => n2181, Z => n254);
   U261 : BUF_X1 port map( A => n2176, Z => n242);
   U262 : BUF_X1 port map( A => n49, Z => n170);
   U263 : BUF_X1 port map( A => n51, Z => n182);
   U264 : BUF_X1 port map( A => n52, Z => n110);
   U265 : BUF_X1 port map( A => n53, Z => n122);
   U266 : BUF_X1 port map( A => n55, Z => n134);
   U267 : BUF_X1 port map( A => n41, Z => n146);
   U268 : BUF_X1 port map( A => n59, Z => n272);
   U269 : BUF_X1 port map( A => n56, Z => n98);
   U270 : BUF_X1 port map( A => n60, Z => n284);
   U271 : BUF_X1 port map( A => n47, Z => n212);
   U272 : BUF_X1 port map( A => n48, Z => n224);
   U273 : BUF_X1 port map( A => n50, Z => n236);
   U274 : BUF_X1 port map( A => n42, Z => n248);
   U275 : BUF_X1 port map( A => n54, Z => n200);
   U276 : BUF_X1 port map( A => n1025, Z => n164);
   U277 : BUF_X1 port map( A => n1028, Z => n176);
   U278 : BUF_X1 port map( A => n1006, Z => n104);
   U279 : BUF_X1 port map( A => n1009, Z => n116);
   U280 : BUF_X1 port map( A => n1003, Z => n92);
   U281 : BUF_X1 port map( A => n1022, Z => n152);
   U282 : BUF_X1 port map( A => n1019, Z => n140);
   U283 : BUF_X1 port map( A => n1026, Z => n167);
   U284 : BUF_X1 port map( A => n1029, Z => n179);
   U285 : BUF_X1 port map( A => n1007, Z => n107);
   U286 : BUF_X1 port map( A => n1010, Z => n119);
   U287 : BUF_X1 port map( A => n1013, Z => n131);
   U288 : BUF_X1 port map( A => n1004, Z => n95);
   U289 : BUF_X1 port map( A => n1023, Z => n155);
   U290 : BUF_X1 port map( A => n1020, Z => n143);
   U291 : BUF_X1 port map( A => n43, Z => n173);
   U292 : BUF_X1 port map( A => n44, Z => n185);
   U293 : BUF_X1 port map( A => n39, Z => n161);
   U294 : BUF_X1 port map( A => n65, Z => n113);
   U295 : BUF_X1 port map( A => n62, Z => n125);
   U296 : BUF_X1 port map( A => n66, Z => n137);
   U297 : BUF_X1 port map( A => n37, Z => n149);
   U298 : BUF_X1 port map( A => n46, Z => n101);
   U299 : BUF_X1 port map( A => n57, Z => n275);
   U300 : BUF_X1 port map( A => n40, Z => n263);
   U301 : BUF_X1 port map( A => n58, Z => n287);
   U302 : BUF_X1 port map( A => n63, Z => n215);
   U303 : BUF_X1 port map( A => n61, Z => n227);
   U304 : BUF_X1 port map( A => n38, Z => n251);
   U305 : BUF_X1 port map( A => n64, Z => n239);
   U306 : BUF_X1 port map( A => n45, Z => n203);
   U307 : AND2_X1 port map( A1 => n85, A2 => n291, ZN => n27);
   U308 : AND2_X1 port map( A1 => n85, A2 => n189, ZN => n28);
   U309 : AND2_X1 port map( A1 => n31, A2 => n33, ZN => n29);
   U310 : AND2_X1 port map( A1 => n32, A2 => n34, ZN => n30);
   U311 : AND2_X2 port map( A1 => n392, A2 => n391, ZN => n31);
   U312 : AND2_X2 port map( A1 => n1044, A2 => n1043, ZN => n32);
   U313 : BUF_X1 port map( A => n1039, Z => n190);
   U314 : BUF_X1 port map( A => n2203, Z => n292);
   U315 : AND2_X1 port map( A1 => n81, A2 => n404, ZN => n33);
   U316 : AND2_X1 port map( A1 => n82, A2 => n1066, ZN => n34);
   U317 : AND3_X1 port map( A1 => n1065, A2 => n1066, A3 => n1048, ZN => n35);
   U318 : AND3_X1 port map( A1 => n403, A2 => n404, A3 => n394, ZN => n36);
   U319 : AND2_X1 port map( A1 => n67, A2 => n69, ZN => n37);
   U320 : AND2_X1 port map( A1 => n68, A2 => n70, ZN => n38);
   U321 : AND2_X1 port map( A1 => n31, A2 => n69, ZN => n39);
   U322 : AND2_X1 port map( A1 => n32, A2 => n70, ZN => n40);
   U323 : AND2_X1 port map( A1 => n33, A2 => n67, ZN => n41);
   U324 : AND2_X1 port map( A1 => n34, A2 => n68, ZN => n42);
   U325 : AND2_X1 port map( A1 => n72, A2 => n1, ZN => n43);
   U326 : AND2_X1 port map( A1 => n72, A2 => n2, ZN => n44);
   U327 : AND2_X1 port map( A1 => n74, A2 => n3, ZN => n45);
   U328 : AND2_X1 port map( A1 => n78, A2 => n1, ZN => n46);
   U329 : AND2_X1 port map( A1 => n75, A2 => n4, ZN => n47);
   U330 : AND2_X1 port map( A1 => n35, A2 => n3, ZN => n48);
   U331 : AND2_X1 port map( A1 => n71, A2 => n1, ZN => n49);
   U332 : AND2_X1 port map( A1 => n35, A2 => n4, ZN => n50);
   U333 : AND2_X1 port map( A1 => n71, A2 => n2, ZN => n51);
   U334 : AND2_X1 port map( A1 => n77, A2 => n2, ZN => n52);
   U335 : AND2_X1 port map( A1 => n36, A2 => n1, ZN => n53);
   U336 : AND2_X1 port map( A1 => n75, A2 => n3, ZN => n54);
   U337 : AND2_X1 port map( A1 => n36, A2 => n2, ZN => n55);
   U338 : AND2_X1 port map( A1 => n77, A2 => n1, ZN => n56);
   U339 : AND2_X1 port map( A1 => n80, A2 => n3, ZN => n57);
   U340 : AND2_X1 port map( A1 => n80, A2 => n4, ZN => n58);
   U341 : AND2_X1 port map( A1 => n79, A2 => n3, ZN => n59);
   U342 : AND2_X1 port map( A1 => n79, A2 => n4, ZN => n60);
   U343 : AND2_X1 port map( A1 => n73, A2 => n3, ZN => n61);
   U344 : AND2_X1 port map( A1 => n76, A2 => n1, ZN => n62);
   U345 : AND2_X1 port map( A1 => n74, A2 => n4, ZN => n63);
   U346 : AND2_X1 port map( A1 => n73, A2 => n4, ZN => n64);
   U347 : AND2_X1 port map( A1 => n78, A2 => n2, ZN => n65);
   U348 : AND2_X1 port map( A1 => n76, A2 => n2, ZN => n66);
   U349 : AND2_X2 port map( A1 => ADD_RD2(2), A2 => n392, ZN => n67);
   U350 : AND2_X2 port map( A1 => ADD_RD1(2), A2 => n1044, ZN => n68);
   U351 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n83, ZN => n4398);
   U352 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n83, ZN => n4400);
   U353 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n83, ZN => n4402);
   U354 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n81, ZN => n69);
   U355 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n82, ZN => n70);
   U356 : AND3_X1 port map( A1 => ADD_RD2(4), A2 => n404, A3 => n403, ZN => n71
                           );
   U357 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n403, ZN 
                           => n72);
   U358 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => n1065, A3 => n1048, ZN => 
                           n73);
   U359 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n1048, ZN
                           => n74);
   U360 : AND3_X1 port map( A1 => ADD_RD1(3), A2 => n1066, A3 => n1048, ZN => 
                           n75);
   U361 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => n403, A3 => n394, ZN => n76
                           );
   U362 : AND3_X1 port map( A1 => ADD_RD2(3), A2 => n404, A3 => n394, ZN => n77
                           );
   U363 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n394, ZN 
                           => n78);
   U364 : AND3_X1 port map( A1 => ADD_RD1(4), A2 => n1066, A3 => n1065, ZN => 
                           n79);
   U365 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n1065, ZN
                           => n80);
   U366 : AND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n81);
   U367 : AND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n82);
   U368 : INV_X1 port map( A => n87, ZN => n83);
   U369 : INV_X1 port map( A => n86, ZN => n84);
   U370 : INV_X1 port map( A => n86, ZN => n85);
   U371 : INV_X1 port map( A => RST, ZN => n86);
   U372 : INV_X1 port map( A => RST, ZN => n87);
   U373 : OR2_X1 port map( A1 => RD2, A2 => n87, ZN => n1039);
   U374 : INV_X1 port map( A => ADD_RD2(4), ZN => n394);
   U375 : INV_X1 port map( A => ADD_RD2(0), ZN => n404);
   U376 : INV_X1 port map( A => ADD_RD2(1), ZN => n392);
   U377 : NAND2_X1 port map( A1 => n78, A2 => n67, ZN => n1004);
   U378 : NAND2_X1 port map( A1 => n77, A2 => n67, ZN => n1003);
   U379 : OAI22_X1 port map( A1 => n1041, A2 => n93, B1 => n1040, B2 => n90, ZN
                           => n390);
   U380 : AOI221_X1 port map( B1 => n99, B2 => n3842, C1 => n96, C2 => n3876, A
                           => n390, ZN => n400);
   U381 : INV_X1 port map( A => ADD_RD2(2), ZN => n391);
   U382 : NAND2_X1 port map( A1 => n78, A2 => n31, ZN => n1007);
   U383 : NAND2_X1 port map( A1 => n77, A2 => n31, ZN => n1006);
   U384 : OAI22_X1 port map( A1 => n1046, A2 => n105, B1 => n1045, B2 => n102, 
                           ZN => n393);
   U385 : AOI221_X1 port map( B1 => n111, B2 => n3978, C1 => n108, C2 => n4012,
                           A => n393, ZN => n399);
   U386 : INV_X1 port map( A => ADD_RD2(3), ZN => n403);
   U387 : NAND2_X1 port map( A1 => n76, A2 => n67, ZN => n1010);
   U388 : NAND2_X1 port map( A1 => n36, A2 => n67, ZN => n1009);
   U389 : OAI22_X1 port map( A1 => n1050, A2 => n117, B1 => n1049, B2 => n114, 
                           ZN => n395);
   U390 : AOI221_X1 port map( B1 => n123, B2 => n4118, C1 => n120, C2 => n4153,
                           A => n395, ZN => n398);
   U391 : NAND2_X1 port map( A1 => n76, A2 => n31, ZN => n1013);
   U392 : NAND2_X1 port map( A1 => n36, A2 => n31, ZN => n1012);
   U393 : OAI22_X1 port map( A1 => n1053, A2 => n129, B1 => n1052, B2 => n126, 
                           ZN => n396);
   U394 : AOI221_X1 port map( B1 => n135, B2 => n4258, C1 => n132, C2 => n4293,
                           A => n396, ZN => n397);
   U395 : NAND4_X1 port map( A1 => n400, A2 => n399, A3 => n398, A4 => n397, ZN
                           => n412);
   U396 : NAND2_X1 port map( A1 => n1, A2 => n69, ZN => n1020);
   U397 : NAND2_X1 port map( A1 => n1, A2 => n33, ZN => n1019);
   U398 : OAI22_X1 port map( A1 => n1060, A2 => n141, B1 => n1059, B2 => n138, 
                           ZN => n401);
   U399 : AOI221_X1 port map( B1 => n147, B2 => n2273, C1 => n144, C2 => n2307,
                           A => n401, ZN => n410);
   U400 : NAND2_X1 port map( A1 => n2, A2 => n69, ZN => n1023);
   U401 : NAND2_X1 port map( A1 => n2, A2 => n33, ZN => n1022);
   U402 : OAI22_X1 port map( A1 => n1063, A2 => n153, B1 => n1062, B2 => n150, 
                           ZN => n402);
   U403 : AOI221_X1 port map( B1 => n159, B2 => n2409, C1 => n156, C2 => n2447,
                           A => n402, ZN => n409);
   U404 : NAND2_X1 port map( A1 => n72, A2 => n67, ZN => n1026);
   U405 : NAND2_X1 port map( A1 => n71, A2 => n67, ZN => n1025);
   U406 : OAI22_X1 port map( A1 => n1068, A2 => n165, B1 => n1067, B2 => n162, 
                           ZN => n405);
   U407 : AOI221_X1 port map( B1 => n171, B2 => n2481, C1 => n168, C2 => n2515,
                           A => n405, ZN => n408);
   U408 : NAND2_X1 port map( A1 => n72, A2 => n31, ZN => n1029);
   U409 : NAND2_X1 port map( A1 => n71, A2 => n31, ZN => n1028);
   U410 : OAI22_X1 port map( A1 => n1071, A2 => n177, B1 => n1070, B2 => n174, 
                           ZN => n406);
   U411 : AOI221_X1 port map( B1 => n183, B2 => n3705, C1 => n180, C2 => n3739,
                           A => n406, ZN => n407);
   U412 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => n411);
   U413 : OAI21_X1 port map( B1 => n412, B2 => n411, A => n186, ZN => n413);
   U414 : OAI21_X1 port map( B1 => n189, B2 => n414, A => n413, ZN => n2527);
   U415 : OAI22_X1 port map( A1 => n1082, A2 => n93, B1 => n1081, B2 => n90, ZN
                           => n415);
   U416 : AOI221_X1 port map( B1 => n99, B2 => n3843, C1 => n96, C2 => n3877, A
                           => n415, ZN => n422);
   U417 : OAI22_X1 port map( A1 => n1085, A2 => n105, B1 => n1084, B2 => n102, 
                           ZN => n416);
   U418 : AOI221_X1 port map( B1 => n111, B2 => n3979, C1 => n108, C2 => n4013,
                           A => n416, ZN => n421);
   U419 : OAI22_X1 port map( A1 => n1088, A2 => n117, B1 => n1087, B2 => n114, 
                           ZN => n417);
   U420 : AOI221_X1 port map( B1 => n123, B2 => n4119, C1 => n120, C2 => n4154,
                           A => n417, ZN => n420);
   U421 : OAI22_X1 port map( A1 => n1091, A2 => n129, B1 => n1090, B2 => n126, 
                           ZN => n418);
   U422 : AOI221_X1 port map( B1 => n135, B2 => n4259, C1 => n132, C2 => n4295,
                           A => n418, ZN => n419);
   U423 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => n432);
   U424 : OAI22_X1 port map( A1 => n1098, A2 => n141, B1 => n1097, B2 => n138, 
                           ZN => n423);
   U425 : AOI221_X1 port map( B1 => n147, B2 => n2274, C1 => n144, C2 => n2308,
                           A => n423, ZN => n430);
   U426 : OAI22_X1 port map( A1 => n1101, A2 => n153, B1 => n1100, B2 => n150, 
                           ZN => n424);
   U427 : AOI221_X1 port map( B1 => n159, B2 => n2410, C1 => n156, C2 => n2448,
                           A => n424, ZN => n429);
   U428 : OAI22_X1 port map( A1 => n1104, A2 => n165, B1 => n1103, B2 => n162, 
                           ZN => n425);
   U429 : AOI221_X1 port map( B1 => n171, B2 => n2482, C1 => n168, C2 => n2516,
                           A => n425, ZN => n428);
   U430 : OAI22_X1 port map( A1 => n1107, A2 => n177, B1 => n1106, B2 => n174, 
                           ZN => n426);
   U431 : AOI221_X1 port map( B1 => n183, B2 => n3706, C1 => n180, C2 => n3740,
                           A => n426, ZN => n427);
   U432 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => n431);
   U433 : OAI21_X1 port map( B1 => n432, B2 => n431, A => n186, ZN => n433);
   U434 : OAI21_X1 port map( B1 => n189, B2 => n89, A => n433, ZN => n2528);
   U435 : OAI22_X1 port map( A1 => n1118, A2 => n93, B1 => n1117, B2 => n90, ZN
                           => n434);
   U436 : AOI221_X1 port map( B1 => n99, B2 => n3844, C1 => n96, C2 => n3878, A
                           => n434, ZN => n441);
   U437 : OAI22_X1 port map( A1 => n1121, A2 => n105, B1 => n1120, B2 => n102, 
                           ZN => n435);
   U438 : AOI221_X1 port map( B1 => n111, B2 => n3980, C1 => n108, C2 => n4014,
                           A => n435, ZN => n440);
   U439 : OAI22_X1 port map( A1 => n1124, A2 => n117, B1 => n1123, B2 => n114, 
                           ZN => n436);
   U440 : AOI221_X1 port map( B1 => n123, B2 => n4120, C1 => n120, C2 => n4155,
                           A => n436, ZN => n439);
   U441 : OAI22_X1 port map( A1 => n1127, A2 => n129, B1 => n1126, B2 => n126, 
                           ZN => n437);
   U442 : AOI221_X1 port map( B1 => n135, B2 => n4260, C1 => n132, C2 => n4297,
                           A => n437, ZN => n438);
   U443 : NAND4_X1 port map( A1 => n441, A2 => n440, A3 => n439, A4 => n438, ZN
                           => n451);
   U444 : OAI22_X1 port map( A1 => n1134, A2 => n141, B1 => n1133, B2 => n138, 
                           ZN => n442);
   U445 : AOI221_X1 port map( B1 => n147, B2 => n2275, C1 => n144, C2 => n2309,
                           A => n442, ZN => n449);
   U446 : OAI22_X1 port map( A1 => n1137, A2 => n153, B1 => n1136, B2 => n150, 
                           ZN => n443);
   U447 : AOI221_X1 port map( B1 => n159, B2 => n2411, C1 => n156, C2 => n2449,
                           A => n443, ZN => n448);
   U448 : OAI22_X1 port map( A1 => n1140, A2 => n165, B1 => n1139, B2 => n162, 
                           ZN => n444);
   U449 : AOI221_X1 port map( B1 => n171, B2 => n2483, C1 => n168, C2 => n2517,
                           A => n444, ZN => n447);
   U450 : OAI22_X1 port map( A1 => n1143, A2 => n177, B1 => n1142, B2 => n174, 
                           ZN => n445);
   U451 : AOI221_X1 port map( B1 => n183, B2 => n3707, C1 => n180, C2 => n3741,
                           A => n445, ZN => n446);
   U452 : NAND4_X1 port map( A1 => n449, A2 => n448, A3 => n447, A4 => n446, ZN
                           => n450);
   U453 : OAI21_X1 port map( B1 => n451, B2 => n450, A => n186, ZN => n452);
   U454 : OAI21_X1 port map( B1 => n189, B2 => n88, A => n452, ZN => n2529);
   U455 : OAI22_X1 port map( A1 => n1154, A2 => n93, B1 => n1153, B2 => n90, ZN
                           => n453);
   U456 : AOI221_X1 port map( B1 => n99, B2 => n3845, C1 => n96, C2 => n3879, A
                           => n453, ZN => n460);
   U457 : OAI22_X1 port map( A1 => n1157, A2 => n105, B1 => n1156, B2 => n102, 
                           ZN => n454);
   U458 : AOI221_X1 port map( B1 => n111, B2 => n3981, C1 => n108, C2 => n4015,
                           A => n454, ZN => n459);
   U459 : OAI22_X1 port map( A1 => n1160, A2 => n117, B1 => n1159, B2 => n114, 
                           ZN => n455);
   U460 : AOI221_X1 port map( B1 => n123, B2 => n4121, C1 => n120, C2 => n4156,
                           A => n455, ZN => n458);
   U461 : OAI22_X1 port map( A1 => n1163, A2 => n129, B1 => n1162, B2 => n126, 
                           ZN => n456);
   U462 : AOI221_X1 port map( B1 => n135, B2 => n4261, C1 => n132, C2 => n4299,
                           A => n456, ZN => n457);
   U463 : NAND4_X1 port map( A1 => n460, A2 => n459, A3 => n458, A4 => n457, ZN
                           => n470);
   U464 : OAI22_X1 port map( A1 => n1170, A2 => n141, B1 => n1169, B2 => n138, 
                           ZN => n461);
   U465 : AOI221_X1 port map( B1 => n147, B2 => n2276, C1 => n144, C2 => n2310,
                           A => n461, ZN => n468);
   U466 : OAI22_X1 port map( A1 => n1173, A2 => n153, B1 => n1172, B2 => n150, 
                           ZN => n462);
   U467 : AOI221_X1 port map( B1 => n159, B2 => n2412, C1 => n156, C2 => n2450,
                           A => n462, ZN => n467);
   U468 : OAI22_X1 port map( A1 => n1176, A2 => n165, B1 => n1175, B2 => n162, 
                           ZN => n463);
   U469 : AOI221_X1 port map( B1 => n171, B2 => n2484, C1 => n168, C2 => n2518,
                           A => n463, ZN => n466);
   U470 : OAI22_X1 port map( A1 => n1179, A2 => n177, B1 => n1178, B2 => n174, 
                           ZN => n464);
   U471 : AOI221_X1 port map( B1 => n183, B2 => n3708, C1 => n180, C2 => n3742,
                           A => n464, ZN => n465);
   U472 : NAND4_X1 port map( A1 => n468, A2 => n467, A3 => n466, A4 => n465, ZN
                           => n469);
   U473 : OAI21_X1 port map( B1 => n470, B2 => n469, A => n186, ZN => n471);
   U474 : OAI21_X1 port map( B1 => n189, B2 => n472, A => n471, ZN => n2530);
   U475 : OAI22_X1 port map( A1 => n1190, A2 => n93, B1 => n1189, B2 => n90, ZN
                           => n473);
   U476 : AOI221_X1 port map( B1 => n99, B2 => n3846, C1 => n96, C2 => n3880, A
                           => n473, ZN => n480);
   U477 : OAI22_X1 port map( A1 => n1193, A2 => n105, B1 => n1192, B2 => n102, 
                           ZN => n474);
   U478 : AOI221_X1 port map( B1 => n111, B2 => n3982, C1 => n108, C2 => n4016,
                           A => n474, ZN => n479);
   U479 : OAI22_X1 port map( A1 => n1196, A2 => n117, B1 => n1195, B2 => n114, 
                           ZN => n475);
   U480 : AOI221_X1 port map( B1 => n123, B2 => n4122, C1 => n120, C2 => n4157,
                           A => n475, ZN => n478);
   U481 : OAI22_X1 port map( A1 => n1199, A2 => n129, B1 => n1198, B2 => n126, 
                           ZN => n476);
   U482 : AOI221_X1 port map( B1 => n135, B2 => n4262, C1 => n132, C2 => n4301,
                           A => n476, ZN => n477);
   U483 : NAND4_X1 port map( A1 => n480, A2 => n479, A3 => n478, A4 => n477, ZN
                           => n490);
   U484 : OAI22_X1 port map( A1 => n1206, A2 => n141, B1 => n1205, B2 => n138, 
                           ZN => n481);
   U485 : AOI221_X1 port map( B1 => n147, B2 => n2277, C1 => n144, C2 => n2311,
                           A => n481, ZN => n488);
   U486 : OAI22_X1 port map( A1 => n1209, A2 => n153, B1 => n1208, B2 => n150, 
                           ZN => n482);
   U487 : AOI221_X1 port map( B1 => n159, B2 => n2413, C1 => n156, C2 => n2451,
                           A => n482, ZN => n487);
   U488 : OAI22_X1 port map( A1 => n1212, A2 => n165, B1 => n1211, B2 => n162, 
                           ZN => n483);
   U489 : AOI221_X1 port map( B1 => n171, B2 => n2485, C1 => n168, C2 => n2519,
                           A => n483, ZN => n486);
   U490 : OAI22_X1 port map( A1 => n1215, A2 => n177, B1 => n1214, B2 => n174, 
                           ZN => n484);
   U491 : AOI221_X1 port map( B1 => n183, B2 => n3709, C1 => n180, C2 => n3743,
                           A => n484, ZN => n485);
   U492 : NAND4_X1 port map( A1 => n488, A2 => n487, A3 => n486, A4 => n485, ZN
                           => n489);
   U493 : OAI21_X1 port map( B1 => n490, B2 => n489, A => n186, ZN => n491);
   U494 : OAI21_X1 port map( B1 => n189, B2 => n492, A => n491, ZN => n2531);
   U495 : OAI22_X1 port map( A1 => n1226, A2 => n93, B1 => n1225, B2 => n90, ZN
                           => n493);
   U496 : AOI221_X1 port map( B1 => n99, B2 => n3847, C1 => n96, C2 => n3881, A
                           => n493, ZN => n500);
   U497 : OAI22_X1 port map( A1 => n1229, A2 => n105, B1 => n1228, B2 => n102, 
                           ZN => n494);
   U498 : AOI221_X1 port map( B1 => n111, B2 => n3983, C1 => n108, C2 => n4017,
                           A => n494, ZN => n499);
   U499 : OAI22_X1 port map( A1 => n1232, A2 => n117, B1 => n1231, B2 => n114, 
                           ZN => n495);
   U500 : AOI221_X1 port map( B1 => n123, B2 => n4123, C1 => n120, C2 => n4158,
                           A => n495, ZN => n498);
   U501 : OAI22_X1 port map( A1 => n1235, A2 => n129, B1 => n1234, B2 => n126, 
                           ZN => n496);
   U502 : AOI221_X1 port map( B1 => n135, B2 => n4263, C1 => n132, C2 => n4303,
                           A => n496, ZN => n497);
   U503 : NAND4_X1 port map( A1 => n500, A2 => n499, A3 => n498, A4 => n497, ZN
                           => n510);
   U504 : OAI22_X1 port map( A1 => n1242, A2 => n141, B1 => n1241, B2 => n138, 
                           ZN => n501);
   U505 : AOI221_X1 port map( B1 => n147, B2 => n2278, C1 => n144, C2 => n2312,
                           A => n501, ZN => n508);
   U506 : OAI22_X1 port map( A1 => n1245, A2 => n153, B1 => n1244, B2 => n150, 
                           ZN => n502);
   U507 : AOI221_X1 port map( B1 => n159, B2 => n2414, C1 => n156, C2 => n2452,
                           A => n502, ZN => n507);
   U508 : OAI22_X1 port map( A1 => n1248, A2 => n165, B1 => n1247, B2 => n162, 
                           ZN => n503);
   U509 : AOI221_X1 port map( B1 => n171, B2 => n2486, C1 => n168, C2 => n2520,
                           A => n503, ZN => n506);
   U510 : OAI22_X1 port map( A1 => n1251, A2 => n177, B1 => n1250, B2 => n174, 
                           ZN => n504);
   U511 : AOI221_X1 port map( B1 => n183, B2 => n3710, C1 => n180, C2 => n3744,
                           A => n504, ZN => n505);
   U512 : NAND4_X1 port map( A1 => n508, A2 => n507, A3 => n506, A4 => n505, ZN
                           => n509);
   U513 : OAI21_X1 port map( B1 => n510, B2 => n509, A => n186, ZN => n511);
   U514 : OAI21_X1 port map( B1 => n189, B2 => n512, A => n511, ZN => n2532);
   U515 : OAI22_X1 port map( A1 => n1262, A2 => n93, B1 => n1261, B2 => n90, ZN
                           => n513);
   U516 : AOI221_X1 port map( B1 => n99, B2 => n3848, C1 => n96, C2 => n3882, A
                           => n513, ZN => n520);
   U517 : OAI22_X1 port map( A1 => n1265, A2 => n105, B1 => n1264, B2 => n102, 
                           ZN => n514);
   U518 : AOI221_X1 port map( B1 => n111, B2 => n3984, C1 => n108, C2 => n4018,
                           A => n514, ZN => n519);
   U519 : OAI22_X1 port map( A1 => n1268, A2 => n117, B1 => n1267, B2 => n114, 
                           ZN => n515);
   U520 : AOI221_X1 port map( B1 => n123, B2 => n4124, C1 => n120, C2 => n4159,
                           A => n515, ZN => n518);
   U521 : OAI22_X1 port map( A1 => n1271, A2 => n129, B1 => n1270, B2 => n126, 
                           ZN => n516);
   U522 : AOI221_X1 port map( B1 => n135, B2 => n4264, C1 => n132, C2 => n4305,
                           A => n516, ZN => n517);
   U523 : NAND4_X1 port map( A1 => n520, A2 => n519, A3 => n518, A4 => n517, ZN
                           => n530);
   U524 : OAI22_X1 port map( A1 => n1278, A2 => n141, B1 => n1277, B2 => n138, 
                           ZN => n521);
   U525 : AOI221_X1 port map( B1 => n147, B2 => n2279, C1 => n144, C2 => n2313,
                           A => n521, ZN => n528);
   U526 : OAI22_X1 port map( A1 => n1281, A2 => n153, B1 => n1280, B2 => n150, 
                           ZN => n522);
   U527 : AOI221_X1 port map( B1 => n159, B2 => n2415, C1 => n156, C2 => n2453,
                           A => n522, ZN => n527);
   U528 : OAI22_X1 port map( A1 => n1284, A2 => n165, B1 => n1283, B2 => n162, 
                           ZN => n523);
   U529 : AOI221_X1 port map( B1 => n171, B2 => n2487, C1 => n168, C2 => n2521,
                           A => n523, ZN => n526);
   U530 : OAI22_X1 port map( A1 => n1287, A2 => n177, B1 => n1286, B2 => n174, 
                           ZN => n524);
   U531 : AOI221_X1 port map( B1 => n183, B2 => n3711, C1 => n180, C2 => n3745,
                           A => n524, ZN => n525);
   U532 : NAND4_X1 port map( A1 => n528, A2 => n527, A3 => n526, A4 => n525, ZN
                           => n529);
   U533 : OAI21_X1 port map( B1 => n530, B2 => n529, A => n186, ZN => n531);
   U534 : OAI21_X1 port map( B1 => n189, B2 => n7, A => n531, ZN => n2533);
   U535 : OAI22_X1 port map( A1 => n1298, A2 => n93, B1 => n1297, B2 => n90, ZN
                           => n532);
   U536 : AOI221_X1 port map( B1 => n99, B2 => n3849, C1 => n96, C2 => n3883, A
                           => n532, ZN => n539);
   U537 : OAI22_X1 port map( A1 => n1301, A2 => n105, B1 => n1300, B2 => n102, 
                           ZN => n533);
   U538 : AOI221_X1 port map( B1 => n111, B2 => n3985, C1 => n108, C2 => n4019,
                           A => n533, ZN => n538);
   U539 : OAI22_X1 port map( A1 => n1304, A2 => n117, B1 => n1303, B2 => n114, 
                           ZN => n534);
   U540 : AOI221_X1 port map( B1 => n123, B2 => n4125, C1 => n120, C2 => n4160,
                           A => n534, ZN => n537);
   U541 : OAI22_X1 port map( A1 => n1307, A2 => n129, B1 => n1306, B2 => n126, 
                           ZN => n535);
   U542 : AOI221_X1 port map( B1 => n135, B2 => n4265, C1 => n132, C2 => n4307,
                           A => n535, ZN => n536);
   U543 : NAND4_X1 port map( A1 => n539, A2 => n538, A3 => n537, A4 => n536, ZN
                           => n549);
   U544 : OAI22_X1 port map( A1 => n1314, A2 => n141, B1 => n1313, B2 => n138, 
                           ZN => n540);
   U545 : AOI221_X1 port map( B1 => n147, B2 => n2280, C1 => n144, C2 => n2314,
                           A => n540, ZN => n547);
   U546 : OAI22_X1 port map( A1 => n1317, A2 => n153, B1 => n1316, B2 => n150, 
                           ZN => n541);
   U547 : AOI221_X1 port map( B1 => n159, B2 => n2416, C1 => n156, C2 => n2454,
                           A => n541, ZN => n546);
   U548 : OAI22_X1 port map( A1 => n1320, A2 => n165, B1 => n1319, B2 => n162, 
                           ZN => n542);
   U549 : AOI221_X1 port map( B1 => n171, B2 => n2488, C1 => n168, C2 => n2522,
                           A => n542, ZN => n545);
   U550 : OAI22_X1 port map( A1 => n1323, A2 => n177, B1 => n1322, B2 => n174, 
                           ZN => n543);
   U551 : AOI221_X1 port map( B1 => n183, B2 => n3712, C1 => n180, C2 => n3746,
                           A => n543, ZN => n544);
   U552 : NAND4_X1 port map( A1 => n547, A2 => n546, A3 => n545, A4 => n544, ZN
                           => n548);
   U553 : OAI21_X1 port map( B1 => n549, B2 => n548, A => n186, ZN => n550);
   U554 : OAI21_X1 port map( B1 => n189, B2 => n8, A => n550, ZN => n2534);
   U555 : OAI22_X1 port map( A1 => n1334, A2 => n93, B1 => n1333, B2 => n90, ZN
                           => n551);
   U556 : AOI221_X1 port map( B1 => n99, B2 => n3850, C1 => n96, C2 => n3884, A
                           => n551, ZN => n558);
   U557 : OAI22_X1 port map( A1 => n1337, A2 => n105, B1 => n1336, B2 => n102, 
                           ZN => n552);
   U558 : AOI221_X1 port map( B1 => n111, B2 => n3986, C1 => n108, C2 => n4020,
                           A => n552, ZN => n557);
   U559 : OAI22_X1 port map( A1 => n1340, A2 => n117, B1 => n1339, B2 => n114, 
                           ZN => n553);
   U560 : AOI221_X1 port map( B1 => n123, B2 => n4126, C1 => n120, C2 => n4161,
                           A => n553, ZN => n556);
   U561 : OAI22_X1 port map( A1 => n1343, A2 => n129, B1 => n1342, B2 => n126, 
                           ZN => n554);
   U562 : AOI221_X1 port map( B1 => n135, B2 => n4266, C1 => n132, C2 => n4309,
                           A => n554, ZN => n555);
   U563 : NAND4_X1 port map( A1 => n558, A2 => n557, A3 => n556, A4 => n555, ZN
                           => n568);
   U564 : OAI22_X1 port map( A1 => n1350, A2 => n141, B1 => n1349, B2 => n138, 
                           ZN => n559);
   U565 : AOI221_X1 port map( B1 => n147, B2 => n2281, C1 => n144, C2 => n2315,
                           A => n559, ZN => n566);
   U566 : OAI22_X1 port map( A1 => n1353, A2 => n153, B1 => n1352, B2 => n150, 
                           ZN => n560);
   U567 : AOI221_X1 port map( B1 => n159, B2 => n2417, C1 => n156, C2 => n2455,
                           A => n560, ZN => n565);
   U568 : OAI22_X1 port map( A1 => n1356, A2 => n165, B1 => n1355, B2 => n162, 
                           ZN => n561);
   U569 : AOI221_X1 port map( B1 => n171, B2 => n2489, C1 => n168, C2 => n2523,
                           A => n561, ZN => n564);
   U570 : OAI22_X1 port map( A1 => n1359, A2 => n177, B1 => n1358, B2 => n174, 
                           ZN => n562);
   U571 : AOI221_X1 port map( B1 => n183, B2 => n3713, C1 => n180, C2 => n3747,
                           A => n562, ZN => n563);
   U572 : NAND4_X1 port map( A1 => n566, A2 => n565, A3 => n564, A4 => n563, ZN
                           => n567);
   U573 : OAI21_X1 port map( B1 => n568, B2 => n567, A => n186, ZN => n569);
   U574 : OAI21_X1 port map( B1 => n189, B2 => n570, A => n569, ZN => n2535);
   U575 : OAI22_X1 port map( A1 => n1369, A2 => n93, B1 => n1368, B2 => n90, ZN
                           => n571);
   U576 : AOI221_X1 port map( B1 => n99, B2 => n3851, C1 => n96, C2 => n3885, A
                           => n571, ZN => n578);
   U577 : OAI22_X1 port map( A1 => n1372, A2 => n105, B1 => n1371, B2 => n102, 
                           ZN => n572);
   U578 : AOI221_X1 port map( B1 => n111, B2 => n3987, C1 => n108, C2 => n4021,
                           A => n572, ZN => n577);
   U579 : OAI22_X1 port map( A1 => n1375, A2 => n117, B1 => n1374, B2 => n114, 
                           ZN => n573);
   U580 : AOI221_X1 port map( B1 => n123, B2 => n4127, C1 => n120, C2 => n4162,
                           A => n573, ZN => n576);
   U581 : OAI22_X1 port map( A1 => n1378, A2 => n129, B1 => n1377, B2 => n126, 
                           ZN => n574);
   U582 : AOI221_X1 port map( B1 => n135, B2 => n4267, C1 => n132, C2 => n4311,
                           A => n574, ZN => n575);
   U583 : NAND4_X1 port map( A1 => n578, A2 => n577, A3 => n576, A4 => n575, ZN
                           => n588);
   U584 : OAI22_X1 port map( A1 => n1385, A2 => n141, B1 => n1384, B2 => n138, 
                           ZN => n579);
   U585 : AOI221_X1 port map( B1 => n147, B2 => n2282, C1 => n144, C2 => n2316,
                           A => n579, ZN => n586);
   U586 : OAI22_X1 port map( A1 => n1388, A2 => n153, B1 => n1387, B2 => n150, 
                           ZN => n580);
   U587 : AOI221_X1 port map( B1 => n159, B2 => n2418, C1 => n156, C2 => n2456,
                           A => n580, ZN => n585);
   U588 : OAI22_X1 port map( A1 => n1391, A2 => n165, B1 => n1390, B2 => n162, 
                           ZN => n581);
   U589 : AOI221_X1 port map( B1 => n171, B2 => n2490, C1 => n168, C2 => n2524,
                           A => n581, ZN => n584);
   U590 : OAI22_X1 port map( A1 => n1394, A2 => n177, B1 => n1393, B2 => n174, 
                           ZN => n582);
   U591 : AOI221_X1 port map( B1 => n183, B2 => n3714, C1 => n180, C2 => n3748,
                           A => n582, ZN => n583);
   U592 : NAND4_X1 port map( A1 => n586, A2 => n585, A3 => n584, A4 => n583, ZN
                           => n587);
   U593 : OAI21_X1 port map( B1 => n588, B2 => n587, A => n186, ZN => n589);
   U594 : OAI21_X1 port map( B1 => n189, B2 => n590, A => n589, ZN => n2536);
   U595 : OAI22_X1 port map( A1 => n1404, A2 => n93, B1 => n1403, B2 => n90, ZN
                           => n591);
   U596 : AOI221_X1 port map( B1 => n99, B2 => n3852, C1 => n96, C2 => n3886, A
                           => n591, ZN => n598);
   U597 : OAI22_X1 port map( A1 => n1407, A2 => n105, B1 => n1406, B2 => n102, 
                           ZN => n592);
   U598 : AOI221_X1 port map( B1 => n111, B2 => n3988, C1 => n108, C2 => n4022,
                           A => n592, ZN => n597);
   U599 : OAI22_X1 port map( A1 => n1410, A2 => n117, B1 => n1409, B2 => n114, 
                           ZN => n593);
   U600 : AOI221_X1 port map( B1 => n123, B2 => n4128, C1 => n120, C2 => n4163,
                           A => n593, ZN => n596);
   U601 : OAI22_X1 port map( A1 => n1413, A2 => n129, B1 => n1412, B2 => n126, 
                           ZN => n594);
   U602 : AOI221_X1 port map( B1 => n135, B2 => n4268, C1 => n132, C2 => n4313,
                           A => n594, ZN => n595);
   U603 : NAND4_X1 port map( A1 => n598, A2 => n597, A3 => n596, A4 => n595, ZN
                           => n608);
   U604 : OAI22_X1 port map( A1 => n1420, A2 => n141, B1 => n1419, B2 => n138, 
                           ZN => n599);
   U605 : AOI221_X1 port map( B1 => n147, B2 => n2283, C1 => n144, C2 => n2317,
                           A => n599, ZN => n606);
   U606 : OAI22_X1 port map( A1 => n1423, A2 => n153, B1 => n1422, B2 => n150, 
                           ZN => n600);
   U607 : AOI221_X1 port map( B1 => n159, B2 => n2419, C1 => n156, C2 => n2457,
                           A => n600, ZN => n605);
   U608 : OAI22_X1 port map( A1 => n1426, A2 => n165, B1 => n1425, B2 => n162, 
                           ZN => n601);
   U609 : AOI221_X1 port map( B1 => n171, B2 => n2491, C1 => n168, C2 => n2525,
                           A => n601, ZN => n604);
   U610 : OAI22_X1 port map( A1 => n1429, A2 => n177, B1 => n1428, B2 => n174, 
                           ZN => n602);
   U611 : AOI221_X1 port map( B1 => n183, B2 => n3715, C1 => n180, C2 => n3749,
                           A => n602, ZN => n603);
   U612 : NAND4_X1 port map( A1 => n606, A2 => n605, A3 => n604, A4 => n603, ZN
                           => n607);
   U613 : OAI21_X1 port map( B1 => n608, B2 => n607, A => n186, ZN => n609);
   U614 : OAI21_X1 port map( B1 => n189, B2 => n20, A => n609, ZN => n2537);
   U615 : OAI22_X1 port map( A1 => n1439, A2 => n93, B1 => n1438, B2 => n90, ZN
                           => n610);
   U616 : AOI221_X1 port map( B1 => n99, B2 => n3853, C1 => n96, C2 => n3887, A
                           => n610, ZN => n617);
   U617 : OAI22_X1 port map( A1 => n1442, A2 => n105, B1 => n1441, B2 => n102, 
                           ZN => n611);
   U618 : AOI221_X1 port map( B1 => n111, B2 => n3989, C1 => n108, C2 => n4023,
                           A => n611, ZN => n616);
   U619 : OAI22_X1 port map( A1 => n1445, A2 => n117, B1 => n1444, B2 => n114, 
                           ZN => n612);
   U620 : AOI221_X1 port map( B1 => n123, B2 => n4129, C1 => n120, C2 => n4164,
                           A => n612, ZN => n615);
   U621 : OAI22_X1 port map( A1 => n1448, A2 => n129, B1 => n1447, B2 => n126, 
                           ZN => n613);
   U622 : AOI221_X1 port map( B1 => n135, B2 => n4269, C1 => n132, C2 => n4315,
                           A => n613, ZN => n614);
   U623 : NAND4_X1 port map( A1 => n617, A2 => n616, A3 => n615, A4 => n614, ZN
                           => n627);
   U624 : OAI22_X1 port map( A1 => n1455, A2 => n141, B1 => n1454, B2 => n138, 
                           ZN => n618);
   U625 : AOI221_X1 port map( B1 => n147, B2 => n2284, C1 => n144, C2 => n2318,
                           A => n618, ZN => n625);
   U626 : OAI22_X1 port map( A1 => n1458, A2 => n153, B1 => n1457, B2 => n150, 
                           ZN => n619);
   U627 : AOI221_X1 port map( B1 => n159, B2 => n2420, C1 => n156, C2 => n2458,
                           A => n619, ZN => n624);
   U628 : OAI22_X1 port map( A1 => n1461, A2 => n165, B1 => n1460, B2 => n162, 
                           ZN => n620);
   U629 : AOI221_X1 port map( B1 => n171, B2 => n2492, C1 => n168, C2 => n2526,
                           A => n620, ZN => n623);
   U630 : OAI22_X1 port map( A1 => n1464, A2 => n177, B1 => n1463, B2 => n174, 
                           ZN => n621);
   U631 : AOI221_X1 port map( B1 => n183, B2 => n3716, C1 => n180, C2 => n3750,
                           A => n621, ZN => n622);
   U632 : NAND4_X1 port map( A1 => n625, A2 => n624, A3 => n623, A4 => n622, ZN
                           => n626);
   U633 : OAI21_X1 port map( B1 => n627, B2 => n626, A => n186, ZN => n628);
   U634 : OAI21_X1 port map( B1 => n190, B2 => n9, A => n628, ZN => n2538);
   U635 : OAI22_X1 port map( A1 => n1474, A2 => n94, B1 => n1473, B2 => n91, ZN
                           => n629);
   U636 : AOI221_X1 port map( B1 => n100, B2 => n3854, C1 => n97, C2 => n3888, 
                           A => n629, ZN => n636);
   U637 : OAI22_X1 port map( A1 => n1477, A2 => n106, B1 => n1476, B2 => n103, 
                           ZN => n630);
   U638 : AOI221_X1 port map( B1 => n112, B2 => n3990, C1 => n109, C2 => n4024,
                           A => n630, ZN => n635);
   U639 : OAI22_X1 port map( A1 => n1480, A2 => n118, B1 => n1479, B2 => n115, 
                           ZN => n631);
   U640 : AOI221_X1 port map( B1 => n124, B2 => n4130, C1 => n121, C2 => n4165,
                           A => n631, ZN => n634);
   U641 : OAI22_X1 port map( A1 => n1483, A2 => n130, B1 => n1482, B2 => n127, 
                           ZN => n632);
   U642 : AOI221_X1 port map( B1 => n136, B2 => n4270, C1 => n133, C2 => n4317,
                           A => n632, ZN => n633);
   U643 : NAND4_X1 port map( A1 => n636, A2 => n635, A3 => n634, A4 => n633, ZN
                           => n646);
   U644 : OAI22_X1 port map( A1 => n1490, A2 => n142, B1 => n1489, B2 => n139, 
                           ZN => n637);
   U645 : AOI221_X1 port map( B1 => n148, B2 => n2285, C1 => n145, C2 => n2319,
                           A => n637, ZN => n644);
   U646 : OAI22_X1 port map( A1 => n1493, A2 => n154, B1 => n1492, B2 => n151, 
                           ZN => n638);
   U647 : AOI221_X1 port map( B1 => n160, B2 => n2421, C1 => n157, C2 => n2459,
                           A => n638, ZN => n643);
   U648 : OAI22_X1 port map( A1 => n1496, A2 => n166, B1 => n1495, B2 => n163, 
                           ZN => n639);
   U649 : AOI221_X1 port map( B1 => n172, B2 => n2493, C1 => n169, C2 => n3615,
                           A => n639, ZN => n642);
   U650 : OAI22_X1 port map( A1 => n1499, A2 => n178, B1 => n1498, B2 => n175, 
                           ZN => n640);
   U651 : AOI221_X1 port map( B1 => n184, B2 => n3717, C1 => n181, C2 => n3751,
                           A => n640, ZN => n641);
   U652 : NAND4_X1 port map( A1 => n644, A2 => n643, A3 => n642, A4 => n641, ZN
                           => n645);
   U653 : OAI21_X1 port map( B1 => n646, B2 => n645, A => n187, ZN => n647);
   U654 : OAI21_X1 port map( B1 => n190, B2 => n648, A => n647, ZN => n2539);
   U655 : OAI22_X1 port map( A1 => n1509, A2 => n94, B1 => n1508, B2 => n91, ZN
                           => n649);
   U656 : AOI221_X1 port map( B1 => n100, B2 => n3855, C1 => n97, C2 => n3889, 
                           A => n649, ZN => n656);
   U657 : OAI22_X1 port map( A1 => n1512, A2 => n106, B1 => n1511, B2 => n103, 
                           ZN => n650);
   U658 : AOI221_X1 port map( B1 => n112, B2 => n3991, C1 => n109, C2 => n4025,
                           A => n650, ZN => n655);
   U659 : OAI22_X1 port map( A1 => n1515, A2 => n118, B1 => n1514, B2 => n115, 
                           ZN => n651);
   U660 : AOI221_X1 port map( B1 => n124, B2 => n4131, C1 => n121, C2 => n4166,
                           A => n651, ZN => n654);
   U661 : OAI22_X1 port map( A1 => n1518, A2 => n130, B1 => n1517, B2 => n127, 
                           ZN => n652);
   U662 : AOI221_X1 port map( B1 => n136, B2 => n4271, C1 => n133, C2 => n4319,
                           A => n652, ZN => n653);
   U663 : NAND4_X1 port map( A1 => n656, A2 => n655, A3 => n654, A4 => n653, ZN
                           => n666);
   U664 : OAI22_X1 port map( A1 => n1525, A2 => n142, B1 => n1524, B2 => n139, 
                           ZN => n657);
   U665 : AOI221_X1 port map( B1 => n148, B2 => n2286, C1 => n145, C2 => n2320,
                           A => n657, ZN => n664);
   U666 : OAI22_X1 port map( A1 => n1528, A2 => n154, B1 => n1527, B2 => n151, 
                           ZN => n658);
   U667 : AOI221_X1 port map( B1 => n160, B2 => n2422, C1 => n157, C2 => n2460,
                           A => n658, ZN => n663);
   U668 : OAI22_X1 port map( A1 => n1531, A2 => n166, B1 => n1530, B2 => n163, 
                           ZN => n659);
   U669 : AOI221_X1 port map( B1 => n172, B2 => n2494, C1 => n169, C2 => n3616,
                           A => n659, ZN => n662);
   U670 : OAI22_X1 port map( A1 => n1534, A2 => n178, B1 => n1533, B2 => n175, 
                           ZN => n660);
   U671 : AOI221_X1 port map( B1 => n184, B2 => n3718, C1 => n181, C2 => n3752,
                           A => n660, ZN => n661);
   U672 : NAND4_X1 port map( A1 => n664, A2 => n663, A3 => n662, A4 => n661, ZN
                           => n665);
   U673 : OAI21_X1 port map( B1 => n666, B2 => n665, A => n187, ZN => n667);
   U674 : OAI21_X1 port map( B1 => n190, B2 => n668, A => n667, ZN => n2540);
   U675 : OAI22_X1 port map( A1 => n1545, A2 => n94, B1 => n1544, B2 => n91, ZN
                           => n669);
   U676 : AOI221_X1 port map( B1 => n100, B2 => n3856, C1 => n97, C2 => n3890, 
                           A => n669, ZN => n676);
   U677 : OAI22_X1 port map( A1 => n1548, A2 => n106, B1 => n1547, B2 => n103, 
                           ZN => n670);
   U678 : AOI221_X1 port map( B1 => n112, B2 => n3992, C1 => n109, C2 => n4026,
                           A => n670, ZN => n675);
   U679 : OAI22_X1 port map( A1 => n1551, A2 => n118, B1 => n1550, B2 => n115, 
                           ZN => n671);
   U680 : AOI221_X1 port map( B1 => n124, B2 => n4132, C1 => n121, C2 => n4167,
                           A => n671, ZN => n674);
   U681 : OAI22_X1 port map( A1 => n1554, A2 => n130, B1 => n1553, B2 => n127, 
                           ZN => n672);
   U682 : AOI221_X1 port map( B1 => n136, B2 => n4272, C1 => n133, C2 => n4321,
                           A => n672, ZN => n673);
   U683 : NAND4_X1 port map( A1 => n676, A2 => n675, A3 => n674, A4 => n673, ZN
                           => n686);
   U684 : OAI22_X1 port map( A1 => n1561, A2 => n142, B1 => n1560, B2 => n139, 
                           ZN => n677);
   U685 : AOI221_X1 port map( B1 => n148, B2 => n2287, C1 => n145, C2 => n2321,
                           A => n677, ZN => n684);
   U686 : OAI22_X1 port map( A1 => n1564, A2 => n154, B1 => n1563, B2 => n151, 
                           ZN => n678);
   U687 : AOI221_X1 port map( B1 => n160, B2 => n2423, C1 => n157, C2 => n2461,
                           A => n678, ZN => n683);
   U688 : OAI22_X1 port map( A1 => n1567, A2 => n166, B1 => n1566, B2 => n163, 
                           ZN => n679);
   U689 : AOI221_X1 port map( B1 => n172, B2 => n2495, C1 => n169, C2 => n3617,
                           A => n679, ZN => n682);
   U690 : OAI22_X1 port map( A1 => n1570, A2 => n178, B1 => n1569, B2 => n175, 
                           ZN => n680);
   U691 : AOI221_X1 port map( B1 => n184, B2 => n3719, C1 => n181, C2 => n3753,
                           A => n680, ZN => n681);
   U692 : NAND4_X1 port map( A1 => n684, A2 => n683, A3 => n682, A4 => n681, ZN
                           => n685);
   U693 : OAI21_X1 port map( B1 => n686, B2 => n685, A => n187, ZN => n687);
   U694 : OAI21_X1 port map( B1 => n190, B2 => n18, A => n687, ZN => n2541);
   U695 : OAI22_X1 port map( A1 => n1580, A2 => n94, B1 => n1579, B2 => n91, ZN
                           => n688);
   U696 : AOI221_X1 port map( B1 => n100, B2 => n3857, C1 => n97, C2 => n3891, 
                           A => n688, ZN => n695);
   U697 : OAI22_X1 port map( A1 => n1583, A2 => n106, B1 => n1582, B2 => n103, 
                           ZN => n689);
   U698 : AOI221_X1 port map( B1 => n112, B2 => n3993, C1 => n109, C2 => n4027,
                           A => n689, ZN => n694);
   U699 : OAI22_X1 port map( A1 => n1586, A2 => n118, B1 => n1585, B2 => n115, 
                           ZN => n690);
   U700 : AOI221_X1 port map( B1 => n124, B2 => n4133, C1 => n121, C2 => n4168,
                           A => n690, ZN => n693);
   U701 : OAI22_X1 port map( A1 => n1589, A2 => n130, B1 => n1588, B2 => n127, 
                           ZN => n691);
   U702 : AOI221_X1 port map( B1 => n136, B2 => n4273, C1 => n133, C2 => n4323,
                           A => n691, ZN => n692);
   U703 : NAND4_X1 port map( A1 => n695, A2 => n694, A3 => n693, A4 => n692, ZN
                           => n705);
   U704 : OAI22_X1 port map( A1 => n1596, A2 => n142, B1 => n1595, B2 => n139, 
                           ZN => n696);
   U705 : AOI221_X1 port map( B1 => n148, B2 => n2288, C1 => n145, C2 => n2322,
                           A => n696, ZN => n703);
   U706 : OAI22_X1 port map( A1 => n1599, A2 => n154, B1 => n1598, B2 => n151, 
                           ZN => n697);
   U707 : AOI221_X1 port map( B1 => n160, B2 => n2424, C1 => n157, C2 => n2462,
                           A => n697, ZN => n702);
   U708 : OAI22_X1 port map( A1 => n1602, A2 => n166, B1 => n1601, B2 => n163, 
                           ZN => n698);
   U709 : AOI221_X1 port map( B1 => n172, B2 => n2496, C1 => n169, C2 => n3618,
                           A => n698, ZN => n701);
   U710 : OAI22_X1 port map( A1 => n1605, A2 => n178, B1 => n1604, B2 => n175, 
                           ZN => n699);
   U711 : AOI221_X1 port map( B1 => n184, B2 => n3720, C1 => n181, C2 => n3754,
                           A => n699, ZN => n700);
   U712 : NAND4_X1 port map( A1 => n703, A2 => n702, A3 => n701, A4 => n700, ZN
                           => n704);
   U713 : OAI21_X1 port map( B1 => n705, B2 => n704, A => n187, ZN => n706);
   U714 : OAI21_X1 port map( B1 => n190, B2 => n707, A => n706, ZN => n2542);
   U715 : OAI22_X1 port map( A1 => n1615, A2 => n94, B1 => n1614, B2 => n91, ZN
                           => n708);
   U716 : AOI221_X1 port map( B1 => n100, B2 => n3858, C1 => n97, C2 => n3892, 
                           A => n708, ZN => n715);
   U717 : OAI22_X1 port map( A1 => n1618, A2 => n106, B1 => n1617, B2 => n103, 
                           ZN => n709);
   U718 : AOI221_X1 port map( B1 => n112, B2 => n3994, C1 => n109, C2 => n4028,
                           A => n709, ZN => n714);
   U719 : OAI22_X1 port map( A1 => n1621, A2 => n118, B1 => n1620, B2 => n115, 
                           ZN => n710);
   U720 : AOI221_X1 port map( B1 => n124, B2 => n4134, C1 => n121, C2 => n4169,
                           A => n710, ZN => n713);
   U721 : OAI22_X1 port map( A1 => n1624, A2 => n130, B1 => n1623, B2 => n127, 
                           ZN => n711);
   U722 : AOI221_X1 port map( B1 => n136, B2 => n4274, C1 => n133, C2 => n4325,
                           A => n711, ZN => n712);
   U723 : NAND4_X1 port map( A1 => n715, A2 => n714, A3 => n713, A4 => n712, ZN
                           => n725);
   U724 : OAI22_X1 port map( A1 => n1631, A2 => n142, B1 => n1630, B2 => n139, 
                           ZN => n716);
   U725 : AOI221_X1 port map( B1 => n148, B2 => n2289, C1 => n145, C2 => n2323,
                           A => n716, ZN => n723);
   U726 : OAI22_X1 port map( A1 => n1634, A2 => n154, B1 => n1633, B2 => n151, 
                           ZN => n717);
   U727 : AOI221_X1 port map( B1 => n160, B2 => n2425, C1 => n157, C2 => n2463,
                           A => n717, ZN => n722);
   U728 : OAI22_X1 port map( A1 => n1637, A2 => n166, B1 => n1636, B2 => n163, 
                           ZN => n718);
   U729 : AOI221_X1 port map( B1 => n172, B2 => n2497, C1 => n169, C2 => n3619,
                           A => n718, ZN => n721);
   U730 : OAI22_X1 port map( A1 => n1640, A2 => n178, B1 => n1639, B2 => n175, 
                           ZN => n719);
   U731 : AOI221_X1 port map( B1 => n184, B2 => n3721, C1 => n181, C2 => n3755,
                           A => n719, ZN => n720);
   U732 : NAND4_X1 port map( A1 => n723, A2 => n722, A3 => n721, A4 => n720, ZN
                           => n724);
   U733 : OAI21_X1 port map( B1 => n725, B2 => n724, A => n187, ZN => n726);
   U734 : OAI21_X1 port map( B1 => n190, B2 => n727, A => n726, ZN => n2543);
   U735 : OAI22_X1 port map( A1 => n1651, A2 => n94, B1 => n1650, B2 => n91, ZN
                           => n728);
   U736 : AOI221_X1 port map( B1 => n100, B2 => n3859, C1 => n97, C2 => n3893, 
                           A => n728, ZN => n735);
   U737 : OAI22_X1 port map( A1 => n1654, A2 => n106, B1 => n1653, B2 => n103, 
                           ZN => n729);
   U738 : AOI221_X1 port map( B1 => n112, B2 => n3995, C1 => n109, C2 => n4029,
                           A => n729, ZN => n734);
   U739 : OAI22_X1 port map( A1 => n1657, A2 => n118, B1 => n1656, B2 => n115, 
                           ZN => n730);
   U740 : AOI221_X1 port map( B1 => n124, B2 => n4135, C1 => n121, C2 => n4170,
                           A => n730, ZN => n733);
   U741 : OAI22_X1 port map( A1 => n1660, A2 => n130, B1 => n1659, B2 => n127, 
                           ZN => n731);
   U742 : AOI221_X1 port map( B1 => n136, B2 => n4275, C1 => n133, C2 => n4327,
                           A => n731, ZN => n732);
   U743 : NAND4_X1 port map( A1 => n735, A2 => n734, A3 => n733, A4 => n732, ZN
                           => n745);
   U744 : OAI22_X1 port map( A1 => n1667, A2 => n142, B1 => n1666, B2 => n139, 
                           ZN => n736);
   U745 : AOI221_X1 port map( B1 => n148, B2 => n2290, C1 => n145, C2 => n2324,
                           A => n736, ZN => n743);
   U746 : OAI22_X1 port map( A1 => n1670, A2 => n154, B1 => n1669, B2 => n151, 
                           ZN => n737);
   U747 : AOI221_X1 port map( B1 => n160, B2 => n2426, C1 => n157, C2 => n2464,
                           A => n737, ZN => n742);
   U748 : OAI22_X1 port map( A1 => n1673, A2 => n166, B1 => n1672, B2 => n163, 
                           ZN => n738);
   U749 : AOI221_X1 port map( B1 => n172, B2 => n2498, C1 => n169, C2 => n3620,
                           A => n738, ZN => n741);
   U750 : OAI22_X1 port map( A1 => n1676, A2 => n178, B1 => n1675, B2 => n175, 
                           ZN => n739);
   U751 : AOI221_X1 port map( B1 => n184, B2 => n3722, C1 => n181, C2 => n3756,
                           A => n739, ZN => n740);
   U752 : NAND4_X1 port map( A1 => n743, A2 => n742, A3 => n741, A4 => n740, ZN
                           => n744);
   U753 : OAI21_X1 port map( B1 => n745, B2 => n744, A => n187, ZN => n746);
   U754 : OAI21_X1 port map( B1 => n190, B2 => n10, A => n746, ZN => n2544);
   U755 : OAI22_X1 port map( A1 => n1687, A2 => n94, B1 => n1686, B2 => n91, ZN
                           => n747);
   U756 : AOI221_X1 port map( B1 => n100, B2 => n3860, C1 => n97, C2 => n3894, 
                           A => n747, ZN => n754);
   U757 : OAI22_X1 port map( A1 => n1690, A2 => n106, B1 => n1689, B2 => n103, 
                           ZN => n748);
   U758 : AOI221_X1 port map( B1 => n112, B2 => n3996, C1 => n109, C2 => n4030,
                           A => n748, ZN => n753);
   U759 : OAI22_X1 port map( A1 => n1693, A2 => n118, B1 => n1692, B2 => n115, 
                           ZN => n749);
   U760 : AOI221_X1 port map( B1 => n124, B2 => n4136, C1 => n121, C2 => n4171,
                           A => n749, ZN => n752);
   U761 : OAI22_X1 port map( A1 => n1696, A2 => n130, B1 => n1695, B2 => n127, 
                           ZN => n750);
   U762 : AOI221_X1 port map( B1 => n136, B2 => n4276, C1 => n133, C2 => n4329,
                           A => n750, ZN => n751);
   U763 : NAND4_X1 port map( A1 => n754, A2 => n753, A3 => n752, A4 => n751, ZN
                           => n764);
   U764 : OAI22_X1 port map( A1 => n1703, A2 => n142, B1 => n1702, B2 => n139, 
                           ZN => n755);
   U765 : AOI221_X1 port map( B1 => n148, B2 => n2291, C1 => n145, C2 => n2325,
                           A => n755, ZN => n762);
   U766 : OAI22_X1 port map( A1 => n1706, A2 => n154, B1 => n1705, B2 => n151, 
                           ZN => n756);
   U767 : AOI221_X1 port map( B1 => n160, B2 => n2427, C1 => n157, C2 => n2465,
                           A => n756, ZN => n761);
   U768 : OAI22_X1 port map( A1 => n1709, A2 => n166, B1 => n1708, B2 => n163, 
                           ZN => n757);
   U769 : AOI221_X1 port map( B1 => n172, B2 => n2499, C1 => n169, C2 => n3621,
                           A => n757, ZN => n760);
   U770 : OAI22_X1 port map( A1 => n1712, A2 => n178, B1 => n1711, B2 => n175, 
                           ZN => n758);
   U771 : AOI221_X1 port map( B1 => n184, B2 => n3723, C1 => n181, C2 => n3757,
                           A => n758, ZN => n759);
   U772 : NAND4_X1 port map( A1 => n762, A2 => n761, A3 => n760, A4 => n759, ZN
                           => n763);
   U773 : OAI21_X1 port map( B1 => n764, B2 => n763, A => n187, ZN => n765);
   U774 : OAI21_X1 port map( B1 => n190, B2 => n11, A => n765, ZN => n2545);
   U775 : OAI22_X1 port map( A1 => n1722, A2 => n94, B1 => n1721, B2 => n91, ZN
                           => n766);
   U776 : AOI221_X1 port map( B1 => n100, B2 => n3861, C1 => n97, C2 => n3895, 
                           A => n766, ZN => n773);
   U777 : OAI22_X1 port map( A1 => n1725, A2 => n106, B1 => n1724, B2 => n103, 
                           ZN => n767);
   U778 : AOI221_X1 port map( B1 => n112, B2 => n3997, C1 => n109, C2 => n4031,
                           A => n767, ZN => n772);
   U779 : OAI22_X1 port map( A1 => n1728, A2 => n118, B1 => n1727, B2 => n115, 
                           ZN => n768);
   U780 : AOI221_X1 port map( B1 => n124, B2 => n4137, C1 => n121, C2 => n4172,
                           A => n768, ZN => n771);
   U781 : OAI22_X1 port map( A1 => n1731, A2 => n130, B1 => n1730, B2 => n127, 
                           ZN => n769);
   U782 : AOI221_X1 port map( B1 => n136, B2 => n4277, C1 => n133, C2 => n4331,
                           A => n769, ZN => n770);
   U783 : NAND4_X1 port map( A1 => n773, A2 => n772, A3 => n771, A4 => n770, ZN
                           => n783);
   U784 : OAI22_X1 port map( A1 => n1738, A2 => n142, B1 => n1737, B2 => n139, 
                           ZN => n774);
   U785 : AOI221_X1 port map( B1 => n148, B2 => n2292, C1 => n145, C2 => n2326,
                           A => n774, ZN => n781);
   U786 : OAI22_X1 port map( A1 => n1741, A2 => n154, B1 => n1740, B2 => n151, 
                           ZN => n775);
   U787 : AOI221_X1 port map( B1 => n160, B2 => n2428, C1 => n157, C2 => n2466,
                           A => n775, ZN => n780);
   U788 : OAI22_X1 port map( A1 => n1744, A2 => n166, B1 => n1743, B2 => n163, 
                           ZN => n776);
   U789 : AOI221_X1 port map( B1 => n172, B2 => n2500, C1 => n169, C2 => n3622,
                           A => n776, ZN => n779);
   U790 : OAI22_X1 port map( A1 => n1747, A2 => n178, B1 => n1746, B2 => n175, 
                           ZN => n777);
   U791 : AOI221_X1 port map( B1 => n184, B2 => n3724, C1 => n181, C2 => n3758,
                           A => n777, ZN => n778);
   U792 : NAND4_X1 port map( A1 => n781, A2 => n780, A3 => n779, A4 => n778, ZN
                           => n782);
   U793 : OAI21_X1 port map( B1 => n783, B2 => n782, A => n187, ZN => n784);
   U794 : OAI21_X1 port map( B1 => n190, B2 => n785, A => n784, ZN => n2546);
   U795 : OAI22_X1 port map( A1 => n1758, A2 => n94, B1 => n1757, B2 => n91, ZN
                           => n786);
   U796 : AOI221_X1 port map( B1 => n100, B2 => n3862, C1 => n97, C2 => n3896, 
                           A => n786, ZN => n793);
   U797 : OAI22_X1 port map( A1 => n1761, A2 => n106, B1 => n1760, B2 => n103, 
                           ZN => n787);
   U798 : AOI221_X1 port map( B1 => n112, B2 => n3998, C1 => n109, C2 => n4032,
                           A => n787, ZN => n792);
   U799 : OAI22_X1 port map( A1 => n1764, A2 => n118, B1 => n1763, B2 => n115, 
                           ZN => n788);
   U800 : AOI221_X1 port map( B1 => n124, B2 => n4138, C1 => n121, C2 => n4173,
                           A => n788, ZN => n791);
   U801 : OAI22_X1 port map( A1 => n1767, A2 => n130, B1 => n1766, B2 => n127, 
                           ZN => n789);
   U802 : AOI221_X1 port map( B1 => n136, B2 => n4278, C1 => n133, C2 => n4333,
                           A => n789, ZN => n790);
   U803 : NAND4_X1 port map( A1 => n793, A2 => n792, A3 => n791, A4 => n790, ZN
                           => n803);
   U804 : OAI22_X1 port map( A1 => n1774, A2 => n142, B1 => n1773, B2 => n139, 
                           ZN => n794);
   U805 : AOI221_X1 port map( B1 => n148, B2 => n2293, C1 => n145, C2 => n2327,
                           A => n794, ZN => n801);
   U806 : OAI22_X1 port map( A1 => n1777, A2 => n154, B1 => n1776, B2 => n151, 
                           ZN => n795);
   U807 : AOI221_X1 port map( B1 => n160, B2 => n2429, C1 => n157, C2 => n2467,
                           A => n795, ZN => n800);
   U808 : OAI22_X1 port map( A1 => n1780, A2 => n166, B1 => n1779, B2 => n163, 
                           ZN => n796);
   U809 : AOI221_X1 port map( B1 => n172, B2 => n2501, C1 => n169, C2 => n3623,
                           A => n796, ZN => n799);
   U810 : OAI22_X1 port map( A1 => n1783, A2 => n178, B1 => n1782, B2 => n175, 
                           ZN => n797);
   U811 : AOI221_X1 port map( B1 => n184, B2 => n3725, C1 => n181, C2 => n3759,
                           A => n797, ZN => n798);
   U812 : NAND4_X1 port map( A1 => n801, A2 => n800, A3 => n799, A4 => n798, ZN
                           => n802);
   U813 : OAI21_X1 port map( B1 => n803, B2 => n802, A => n187, ZN => n804);
   U814 : OAI21_X1 port map( B1 => n190, B2 => n805, A => n804, ZN => n2547);
   U815 : OAI22_X1 port map( A1 => n1794, A2 => n94, B1 => n1793, B2 => n91, ZN
                           => n806);
   U816 : AOI221_X1 port map( B1 => n100, B2 => n3863, C1 => n97, C2 => n3897, 
                           A => n806, ZN => n813);
   U817 : OAI22_X1 port map( A1 => n1797, A2 => n106, B1 => n1796, B2 => n103, 
                           ZN => n807);
   U818 : AOI221_X1 port map( B1 => n112, B2 => n3999, C1 => n109, C2 => n4033,
                           A => n807, ZN => n812);
   U819 : OAI22_X1 port map( A1 => n1800, A2 => n118, B1 => n1799, B2 => n115, 
                           ZN => n808);
   U820 : AOI221_X1 port map( B1 => n124, B2 => n4139, C1 => n121, C2 => n4174,
                           A => n808, ZN => n811);
   U821 : OAI22_X1 port map( A1 => n1803, A2 => n130, B1 => n1802, B2 => n127, 
                           ZN => n809);
   U822 : AOI221_X1 port map( B1 => n136, B2 => n4279, C1 => n133, C2 => n4335,
                           A => n809, ZN => n810);
   U823 : NAND4_X1 port map( A1 => n813, A2 => n812, A3 => n811, A4 => n810, ZN
                           => n823);
   U824 : OAI22_X1 port map( A1 => n1810, A2 => n142, B1 => n1809, B2 => n139, 
                           ZN => n814);
   U825 : AOI221_X1 port map( B1 => n148, B2 => n2294, C1 => n145, C2 => n2328,
                           A => n814, ZN => n821);
   U826 : OAI22_X1 port map( A1 => n1813, A2 => n154, B1 => n1812, B2 => n151, 
                           ZN => n815);
   U827 : AOI221_X1 port map( B1 => n160, B2 => n2430, C1 => n157, C2 => n2468,
                           A => n815, ZN => n820);
   U828 : OAI22_X1 port map( A1 => n1816, A2 => n166, B1 => n1815, B2 => n163, 
                           ZN => n816);
   U829 : AOI221_X1 port map( B1 => n172, B2 => n2502, C1 => n169, C2 => n3624,
                           A => n816, ZN => n819);
   U830 : OAI22_X1 port map( A1 => n1819, A2 => n178, B1 => n1818, B2 => n175, 
                           ZN => n817);
   U831 : AOI221_X1 port map( B1 => n184, B2 => n3726, C1 => n181, C2 => n3760,
                           A => n817, ZN => n818);
   U832 : NAND4_X1 port map( A1 => n821, A2 => n820, A3 => n819, A4 => n818, ZN
                           => n822);
   U833 : OAI21_X1 port map( B1 => n823, B2 => n822, A => n187, ZN => n824);
   U834 : OAI21_X1 port map( B1 => n190, B2 => n13, A => n824, ZN => n2548);
   U835 : OAI22_X1 port map( A1 => n1830, A2 => n94, B1 => n1829, B2 => n91, ZN
                           => n825);
   U836 : AOI221_X1 port map( B1 => n100, B2 => n3864, C1 => n97, C2 => n3898, 
                           A => n825, ZN => n832);
   U837 : OAI22_X1 port map( A1 => n1833, A2 => n106, B1 => n1832, B2 => n103, 
                           ZN => n826);
   U838 : AOI221_X1 port map( B1 => n112, B2 => n4000, C1 => n109, C2 => n4034,
                           A => n826, ZN => n831);
   U839 : OAI22_X1 port map( A1 => n1836, A2 => n118, B1 => n1835, B2 => n115, 
                           ZN => n827);
   U840 : AOI221_X1 port map( B1 => n124, B2 => n4140, C1 => n121, C2 => n4175,
                           A => n827, ZN => n830);
   U841 : OAI22_X1 port map( A1 => n1839, A2 => n130, B1 => n1838, B2 => n127, 
                           ZN => n828);
   U842 : AOI221_X1 port map( B1 => n136, B2 => n4280, C1 => n133, C2 => n4337,
                           A => n828, ZN => n829);
   U843 : NAND4_X1 port map( A1 => n832, A2 => n831, A3 => n830, A4 => n829, ZN
                           => n842);
   U844 : OAI22_X1 port map( A1 => n1846, A2 => n142, B1 => n1845, B2 => n139, 
                           ZN => n833);
   U845 : AOI221_X1 port map( B1 => n148, B2 => n2295, C1 => n145, C2 => n2329,
                           A => n833, ZN => n840);
   U846 : OAI22_X1 port map( A1 => n1849, A2 => n154, B1 => n1848, B2 => n151, 
                           ZN => n834);
   U847 : AOI221_X1 port map( B1 => n160, B2 => n2431, C1 => n157, C2 => n2469,
                           A => n834, ZN => n839);
   U848 : OAI22_X1 port map( A1 => n1852, A2 => n166, B1 => n1851, B2 => n163, 
                           ZN => n835);
   U849 : AOI221_X1 port map( B1 => n172, B2 => n2503, C1 => n169, C2 => n3625,
                           A => n835, ZN => n838);
   U850 : OAI22_X1 port map( A1 => n1855, A2 => n178, B1 => n1854, B2 => n175, 
                           ZN => n836);
   U851 : AOI221_X1 port map( B1 => n184, B2 => n3727, C1 => n181, C2 => n3761,
                           A => n836, ZN => n837);
   U852 : NAND4_X1 port map( A1 => n840, A2 => n839, A3 => n838, A4 => n837, ZN
                           => n841);
   U853 : OAI21_X1 port map( B1 => n842, B2 => n841, A => n187, ZN => n843);
   U854 : OAI21_X1 port map( B1 => n190, B2 => n844, A => n843, ZN => n2549);
   U855 : OAI22_X1 port map( A1 => n1866, A2 => n94, B1 => n1865, B2 => n91, ZN
                           => n845);
   U856 : AOI221_X1 port map( B1 => n100, B2 => n3865, C1 => n97, C2 => n3899, 
                           A => n845, ZN => n852);
   U857 : OAI22_X1 port map( A1 => n1869, A2 => n106, B1 => n1868, B2 => n103, 
                           ZN => n846);
   U858 : AOI221_X1 port map( B1 => n112, B2 => n4001, C1 => n109, C2 => n4035,
                           A => n846, ZN => n851);
   U859 : OAI22_X1 port map( A1 => n1872, A2 => n118, B1 => n1871, B2 => n115, 
                           ZN => n847);
   U860 : AOI221_X1 port map( B1 => n124, B2 => n4141, C1 => n121, C2 => n4176,
                           A => n847, ZN => n850);
   U861 : OAI22_X1 port map( A1 => n1875, A2 => n130, B1 => n1874, B2 => n127, 
                           ZN => n848);
   U862 : AOI221_X1 port map( B1 => n136, B2 => n4281, C1 => n133, C2 => n4339,
                           A => n848, ZN => n849);
   U863 : NAND4_X1 port map( A1 => n852, A2 => n851, A3 => n850, A4 => n849, ZN
                           => n862);
   U864 : OAI22_X1 port map( A1 => n1882, A2 => n142, B1 => n1881, B2 => n139, 
                           ZN => n853);
   U865 : AOI221_X1 port map( B1 => n148, B2 => n2296, C1 => n145, C2 => n2330,
                           A => n853, ZN => n860);
   U866 : OAI22_X1 port map( A1 => n1885, A2 => n154, B1 => n1884, B2 => n151, 
                           ZN => n854);
   U867 : AOI221_X1 port map( B1 => n160, B2 => n2432, C1 => n157, C2 => n2470,
                           A => n854, ZN => n859);
   U868 : OAI22_X1 port map( A1 => n1888, A2 => n166, B1 => n1887, B2 => n163, 
                           ZN => n855);
   U869 : AOI221_X1 port map( B1 => n172, B2 => n2504, C1 => n169, C2 => n3626,
                           A => n855, ZN => n858);
   U870 : OAI22_X1 port map( A1 => n1891, A2 => n178, B1 => n1890, B2 => n175, 
                           ZN => n856);
   U871 : AOI221_X1 port map( B1 => n184, B2 => n3728, C1 => n181, C2 => n3762,
                           A => n856, ZN => n857);
   U872 : NAND4_X1 port map( A1 => n860, A2 => n859, A3 => n858, A4 => n857, ZN
                           => n861);
   U873 : OAI21_X1 port map( B1 => n862, B2 => n861, A => n187, ZN => n863);
   U874 : OAI21_X1 port map( B1 => n191, B2 => n864, A => n863, ZN => n2550);
   U875 : OAI22_X1 port map( A1 => n1902, A2 => n95, B1 => n1901, B2 => n92, ZN
                           => n865);
   U876 : AOI221_X1 port map( B1 => n101, B2 => n3866, C1 => n98, C2 => n3900, 
                           A => n865, ZN => n872);
   U877 : OAI22_X1 port map( A1 => n1905, A2 => n107, B1 => n1904, B2 => n104, 
                           ZN => n866);
   U878 : AOI221_X1 port map( B1 => n113, B2 => n4002, C1 => n110, C2 => n4036,
                           A => n866, ZN => n871);
   U879 : OAI22_X1 port map( A1 => n1908, A2 => n119, B1 => n1907, B2 => n116, 
                           ZN => n867);
   U880 : AOI221_X1 port map( B1 => n125, B2 => n4142, C1 => n122, C2 => n4177,
                           A => n867, ZN => n870);
   U881 : OAI22_X1 port map( A1 => n1911, A2 => n131, B1 => n1910, B2 => n128, 
                           ZN => n868);
   U882 : AOI221_X1 port map( B1 => n137, B2 => n4282, C1 => n134, C2 => n4341,
                           A => n868, ZN => n869);
   U883 : NAND4_X1 port map( A1 => n872, A2 => n871, A3 => n870, A4 => n869, ZN
                           => n882);
   U884 : OAI22_X1 port map( A1 => n1918, A2 => n143, B1 => n1917, B2 => n140, 
                           ZN => n873);
   U885 : AOI221_X1 port map( B1 => n149, B2 => n2297, C1 => n146, C2 => n2331,
                           A => n873, ZN => n880);
   U886 : OAI22_X1 port map( A1 => n1921, A2 => n155, B1 => n1920, B2 => n152, 
                           ZN => n874);
   U887 : AOI221_X1 port map( B1 => n161, B2 => n2433, C1 => n158, C2 => n2471,
                           A => n874, ZN => n879);
   U888 : OAI22_X1 port map( A1 => n1924, A2 => n167, B1 => n1923, B2 => n164, 
                           ZN => n875);
   U889 : AOI221_X1 port map( B1 => n173, B2 => n2505, C1 => n170, C2 => n3627,
                           A => n875, ZN => n878);
   U890 : OAI22_X1 port map( A1 => n1927, A2 => n179, B1 => n1926, B2 => n176, 
                           ZN => n876);
   U891 : AOI221_X1 port map( B1 => n185, B2 => n3729, C1 => n182, C2 => n3763,
                           A => n876, ZN => n877);
   U892 : NAND4_X1 port map( A1 => n880, A2 => n879, A3 => n878, A4 => n877, ZN
                           => n881);
   U893 : OAI21_X1 port map( B1 => n882, B2 => n881, A => n188, ZN => n883);
   U894 : OAI21_X1 port map( B1 => n191, B2 => n14, A => n883, ZN => n2551);
   U895 : OAI22_X1 port map( A1 => n1938, A2 => n95, B1 => n1937, B2 => n92, ZN
                           => n884);
   U896 : AOI221_X1 port map( B1 => n101, B2 => n3867, C1 => n98, C2 => n3901, 
                           A => n884, ZN => n891);
   U897 : OAI22_X1 port map( A1 => n1941, A2 => n107, B1 => n1940, B2 => n104, 
                           ZN => n885);
   U898 : AOI221_X1 port map( B1 => n113, B2 => n4003, C1 => n110, C2 => n4037,
                           A => n885, ZN => n890);
   U899 : OAI22_X1 port map( A1 => n1944, A2 => n119, B1 => n1943, B2 => n116, 
                           ZN => n886);
   U900 : AOI221_X1 port map( B1 => n125, B2 => n4143, C1 => n122, C2 => n4178,
                           A => n886, ZN => n889);
   U901 : OAI22_X1 port map( A1 => n1947, A2 => n131, B1 => n1946, B2 => n128, 
                           ZN => n887);
   U902 : AOI221_X1 port map( B1 => n137, B2 => n4283, C1 => n134, C2 => n4343,
                           A => n887, ZN => n888);
   U903 : NAND4_X1 port map( A1 => n891, A2 => n890, A3 => n889, A4 => n888, ZN
                           => n901);
   U904 : OAI22_X1 port map( A1 => n1954, A2 => n143, B1 => n1953, B2 => n140, 
                           ZN => n892);
   U905 : AOI221_X1 port map( B1 => n149, B2 => n2298, C1 => n146, C2 => n2332,
                           A => n892, ZN => n899);
   U906 : OAI22_X1 port map( A1 => n1957, A2 => n155, B1 => n1956, B2 => n152, 
                           ZN => n893);
   U907 : AOI221_X1 port map( B1 => n161, B2 => n2434, C1 => n158, C2 => n2472,
                           A => n893, ZN => n898);
   U908 : OAI22_X1 port map( A1 => n1960, A2 => n167, B1 => n1959, B2 => n164, 
                           ZN => n894);
   U909 : AOI221_X1 port map( B1 => n173, B2 => n2506, C1 => n170, C2 => n3628,
                           A => n894, ZN => n897);
   U910 : OAI22_X1 port map( A1 => n1963, A2 => n179, B1 => n1962, B2 => n176, 
                           ZN => n895);
   U911 : AOI221_X1 port map( B1 => n185, B2 => n3730, C1 => n182, C2 => n3764,
                           A => n895, ZN => n896);
   U912 : NAND4_X1 port map( A1 => n899, A2 => n898, A3 => n897, A4 => n896, ZN
                           => n900);
   U913 : OAI21_X1 port map( B1 => n901, B2 => n900, A => n188, ZN => n902);
   U914 : OAI21_X1 port map( B1 => n191, B2 => n903, A => n902, ZN => n2552);
   U915 : OAI22_X1 port map( A1 => n1973, A2 => n95, B1 => n1972, B2 => n92, ZN
                           => n904);
   U916 : AOI221_X1 port map( B1 => n101, B2 => n3868, C1 => n98, C2 => n3902, 
                           A => n904, ZN => n911);
   U917 : OAI22_X1 port map( A1 => n1976, A2 => n107, B1 => n1975, B2 => n104, 
                           ZN => n905);
   U918 : AOI221_X1 port map( B1 => n113, B2 => n4004, C1 => n110, C2 => n4038,
                           A => n905, ZN => n910);
   U919 : OAI22_X1 port map( A1 => n1979, A2 => n119, B1 => n1978, B2 => n116, 
                           ZN => n906);
   U920 : AOI221_X1 port map( B1 => n125, B2 => n4144, C1 => n122, C2 => n4179,
                           A => n906, ZN => n909);
   U921 : OAI22_X1 port map( A1 => n1982, A2 => n131, B1 => n1981, B2 => n128, 
                           ZN => n907);
   U922 : AOI221_X1 port map( B1 => n137, B2 => n4284, C1 => n134, C2 => n4345,
                           A => n907, ZN => n908);
   U923 : NAND4_X1 port map( A1 => n911, A2 => n910, A3 => n909, A4 => n908, ZN
                           => n921);
   U924 : OAI22_X1 port map( A1 => n1989, A2 => n143, B1 => n1988, B2 => n140, 
                           ZN => n912);
   U925 : AOI221_X1 port map( B1 => n149, B2 => n2299, C1 => n146, C2 => n2333,
                           A => n912, ZN => n919);
   U926 : OAI22_X1 port map( A1 => n1992, A2 => n155, B1 => n1991, B2 => n152, 
                           ZN => n913);
   U927 : AOI221_X1 port map( B1 => n161, B2 => n2435, C1 => n158, C2 => n2473,
                           A => n913, ZN => n918);
   U928 : OAI22_X1 port map( A1 => n1995, A2 => n167, B1 => n1994, B2 => n164, 
                           ZN => n914);
   U929 : AOI221_X1 port map( B1 => n173, B2 => n2507, C1 => n170, C2 => n3629,
                           A => n914, ZN => n917);
   U930 : OAI22_X1 port map( A1 => n1998, A2 => n179, B1 => n1997, B2 => n176, 
                           ZN => n915);
   U931 : AOI221_X1 port map( B1 => n185, B2 => n3731, C1 => n182, C2 => n3765,
                           A => n915, ZN => n916);
   U932 : NAND4_X1 port map( A1 => n919, A2 => n918, A3 => n917, A4 => n916, ZN
                           => n920);
   U933 : OAI21_X1 port map( B1 => n921, B2 => n920, A => n188, ZN => n922);
   U934 : OAI21_X1 port map( B1 => n191, B2 => n12, A => n922, ZN => n2553);
   U935 : OAI22_X1 port map( A1 => n2008, A2 => n95, B1 => n2007, B2 => n92, ZN
                           => n923);
   U936 : AOI221_X1 port map( B1 => n101, B2 => n3869, C1 => n98, C2 => n3903, 
                           A => n923, ZN => n930);
   U937 : OAI22_X1 port map( A1 => n2011, A2 => n107, B1 => n2010, B2 => n104, 
                           ZN => n924);
   U938 : AOI221_X1 port map( B1 => n113, B2 => n4005, C1 => n110, C2 => n4039,
                           A => n924, ZN => n929);
   U939 : OAI22_X1 port map( A1 => n2014, A2 => n119, B1 => n2013, B2 => n116, 
                           ZN => n925);
   U940 : AOI221_X1 port map( B1 => n125, B2 => n4145, C1 => n122, C2 => n4180,
                           A => n925, ZN => n928);
   U941 : OAI22_X1 port map( A1 => n2017, A2 => n131, B1 => n2016, B2 => n128, 
                           ZN => n926);
   U942 : AOI221_X1 port map( B1 => n137, B2 => n4285, C1 => n134, C2 => n4347,
                           A => n926, ZN => n927);
   U943 : NAND4_X1 port map( A1 => n930, A2 => n929, A3 => n928, A4 => n927, ZN
                           => n940);
   U944 : OAI22_X1 port map( A1 => n2024, A2 => n143, B1 => n2023, B2 => n140, 
                           ZN => n931);
   U945 : AOI221_X1 port map( B1 => n149, B2 => n2300, C1 => n146, C2 => n2334,
                           A => n931, ZN => n938);
   U946 : OAI22_X1 port map( A1 => n2027, A2 => n155, B1 => n2026, B2 => n152, 
                           ZN => n932);
   U947 : AOI221_X1 port map( B1 => n161, B2 => n2436, C1 => n158, C2 => n2474,
                           A => n932, ZN => n937);
   U948 : OAI22_X1 port map( A1 => n2030, A2 => n167, B1 => n2029, B2 => n164, 
                           ZN => n933);
   U949 : AOI221_X1 port map( B1 => n173, B2 => n2508, C1 => n170, C2 => n3630,
                           A => n933, ZN => n936);
   U950 : OAI22_X1 port map( A1 => n2033, A2 => n179, B1 => n2032, B2 => n176, 
                           ZN => n934);
   U951 : AOI221_X1 port map( B1 => n185, B2 => n3732, C1 => n182, C2 => n3766,
                           A => n934, ZN => n935);
   U952 : NAND4_X1 port map( A1 => n938, A2 => n937, A3 => n936, A4 => n935, ZN
                           => n939);
   U953 : OAI21_X1 port map( B1 => n940, B2 => n939, A => n188, ZN => n941);
   U954 : OAI21_X1 port map( B1 => n191, B2 => n942, A => n941, ZN => n2554);
   U955 : OAI22_X1 port map( A1 => n2044, A2 => n95, B1 => n2043, B2 => n92, ZN
                           => n943);
   U956 : AOI221_X1 port map( B1 => n101, B2 => n3870, C1 => n98, C2 => n3904, 
                           A => n943, ZN => n950);
   U957 : OAI22_X1 port map( A1 => n2047, A2 => n107, B1 => n2046, B2 => n104, 
                           ZN => n944);
   U958 : AOI221_X1 port map( B1 => n113, B2 => n4006, C1 => n110, C2 => n4040,
                           A => n944, ZN => n949);
   U959 : OAI22_X1 port map( A1 => n2050, A2 => n119, B1 => n2049, B2 => n116, 
                           ZN => n945);
   U960 : AOI221_X1 port map( B1 => n125, B2 => n4146, C1 => n122, C2 => n4181,
                           A => n945, ZN => n948);
   U961 : OAI22_X1 port map( A1 => n2053, A2 => n131, B1 => n2052, B2 => n128, 
                           ZN => n946);
   U962 : AOI221_X1 port map( B1 => n137, B2 => n4286, C1 => n134, C2 => n4349,
                           A => n946, ZN => n947);
   U963 : NAND4_X1 port map( A1 => n950, A2 => n949, A3 => n948, A4 => n947, ZN
                           => n960);
   U964 : OAI22_X1 port map( A1 => n2060, A2 => n143, B1 => n2059, B2 => n140, 
                           ZN => n951);
   U965 : AOI221_X1 port map( B1 => n149, B2 => n2301, C1 => n146, C2 => n2335,
                           A => n951, ZN => n958);
   U966 : OAI22_X1 port map( A1 => n2063, A2 => n155, B1 => n2062, B2 => n152, 
                           ZN => n952);
   U967 : AOI221_X1 port map( B1 => n161, B2 => n2437, C1 => n158, C2 => n2475,
                           A => n952, ZN => n957);
   U968 : OAI22_X1 port map( A1 => n2066, A2 => n167, B1 => n2065, B2 => n164, 
                           ZN => n953);
   U969 : AOI221_X1 port map( B1 => n173, B2 => n2509, C1 => n170, C2 => n3631,
                           A => n953, ZN => n956);
   U970 : OAI22_X1 port map( A1 => n2069, A2 => n179, B1 => n2068, B2 => n176, 
                           ZN => n954);
   U971 : AOI221_X1 port map( B1 => n185, B2 => n3733, C1 => n182, C2 => n3767,
                           A => n954, ZN => n955);
   U972 : NAND4_X1 port map( A1 => n958, A2 => n957, A3 => n956, A4 => n955, ZN
                           => n959);
   U973 : OAI21_X1 port map( B1 => n960, B2 => n959, A => n188, ZN => n961);
   U974 : OAI21_X1 port map( B1 => n191, B2 => n962, A => n961, ZN => n2555);
   U975 : OAI22_X1 port map( A1 => n2080, A2 => n95, B1 => n2079, B2 => n92, ZN
                           => n963);
   U976 : AOI221_X1 port map( B1 => n101, B2 => n3871, C1 => n98, C2 => n3905, 
                           A => n963, ZN => n970);
   U977 : OAI22_X1 port map( A1 => n2083, A2 => n107, B1 => n2082, B2 => n104, 
                           ZN => n964);
   U978 : AOI221_X1 port map( B1 => n113, B2 => n4007, C1 => n110, C2 => n4041,
                           A => n964, ZN => n969);
   U979 : OAI22_X1 port map( A1 => n2086, A2 => n119, B1 => n2085, B2 => n116, 
                           ZN => n965);
   U980 : AOI221_X1 port map( B1 => n125, B2 => n4147, C1 => n122, C2 => n4182,
                           A => n965, ZN => n968);
   U981 : OAI22_X1 port map( A1 => n2089, A2 => n131, B1 => n2088, B2 => n128, 
                           ZN => n966);
   U982 : AOI221_X1 port map( B1 => n137, B2 => n4287, C1 => n134, C2 => n4351,
                           A => n966, ZN => n967);
   U983 : NAND4_X1 port map( A1 => n970, A2 => n969, A3 => n968, A4 => n967, ZN
                           => n980);
   U984 : OAI22_X1 port map( A1 => n2096, A2 => n143, B1 => n2095, B2 => n140, 
                           ZN => n971);
   U985 : AOI221_X1 port map( B1 => n149, B2 => n2302, C1 => n146, C2 => n2336,
                           A => n971, ZN => n978);
   U986 : OAI22_X1 port map( A1 => n2099, A2 => n155, B1 => n2098, B2 => n152, 
                           ZN => n972);
   U987 : AOI221_X1 port map( B1 => n161, B2 => n2438, C1 => n158, C2 => n2476,
                           A => n972, ZN => n977);
   U988 : OAI22_X1 port map( A1 => n2102, A2 => n167, B1 => n2101, B2 => n164, 
                           ZN => n973);
   U989 : AOI221_X1 port map( B1 => n173, B2 => n2510, C1 => n170, C2 => n3632,
                           A => n973, ZN => n976);
   U990 : OAI22_X1 port map( A1 => n2105, A2 => n179, B1 => n2104, B2 => n176, 
                           ZN => n974);
   U991 : AOI221_X1 port map( B1 => n185, B2 => n3734, C1 => n182, C2 => n3768,
                           A => n974, ZN => n975);
   U992 : NAND4_X1 port map( A1 => n978, A2 => n977, A3 => n976, A4 => n975, ZN
                           => n979);
   U993 : OAI21_X1 port map( B1 => n980, B2 => n979, A => n188, ZN => n981);
   U994 : OAI21_X1 port map( B1 => n191, B2 => n982, A => n981, ZN => n2556);
   U995 : OAI22_X1 port map( A1 => n2116, A2 => n95, B1 => n2115, B2 => n92, ZN
                           => n983);
   U996 : AOI221_X1 port map( B1 => n101, B2 => n3872, C1 => n98, C2 => n3906, 
                           A => n983, ZN => n990);
   U997 : OAI22_X1 port map( A1 => n2119, A2 => n107, B1 => n2118, B2 => n104, 
                           ZN => n984);
   U998 : AOI221_X1 port map( B1 => n113, B2 => n4008, C1 => n110, C2 => n4042,
                           A => n984, ZN => n989);
   U999 : OAI22_X1 port map( A1 => n2122, A2 => n119, B1 => n2121, B2 => n116, 
                           ZN => n985);
   U1000 : AOI221_X1 port map( B1 => n125, B2 => n4148, C1 => n122, C2 => n4183
                           , A => n985, ZN => n988);
   U1001 : OAI22_X1 port map( A1 => n2125, A2 => n131, B1 => n2124, B2 => n128,
                           ZN => n986);
   U1002 : AOI221_X1 port map( B1 => n137, B2 => n4288, C1 => n134, C2 => n4353
                           , A => n986, ZN => n987);
   U1003 : NAND4_X1 port map( A1 => n990, A2 => n989, A3 => n988, A4 => n987, 
                           ZN => n1000);
   U1004 : OAI22_X1 port map( A1 => n2132, A2 => n143, B1 => n2131, B2 => n140,
                           ZN => n991);
   U1005 : AOI221_X1 port map( B1 => n149, B2 => n2303, C1 => n146, C2 => n2337
                           , A => n991, ZN => n998);
   U1006 : OAI22_X1 port map( A1 => n2135, A2 => n155, B1 => n2134, B2 => n152,
                           ZN => n992);
   U1007 : AOI221_X1 port map( B1 => n161, B2 => n2439, C1 => n158, C2 => n2477
                           , A => n992, ZN => n997);
   U1008 : OAI22_X1 port map( A1 => n2138, A2 => n167, B1 => n2137, B2 => n164,
                           ZN => n993);
   U1009 : AOI221_X1 port map( B1 => n173, B2 => n2511, C1 => n170, C2 => n3633
                           , A => n993, ZN => n996);
   U1010 : OAI22_X1 port map( A1 => n2141, A2 => n179, B1 => n2140, B2 => n176,
                           ZN => n994);
   U1011 : AOI221_X1 port map( B1 => n185, B2 => n3735, C1 => n182, C2 => n3769
                           , A => n994, ZN => n995);
   U1012 : NAND4_X1 port map( A1 => n998, A2 => n997, A3 => n996, A4 => n995, 
                           ZN => n999);
   U1013 : OAI21_X1 port map( B1 => n1000, B2 => n999, A => n188, ZN => n1001);
   U1014 : OAI21_X1 port map( B1 => n191, B2 => n1002, A => n1001, ZN => n2557)
                           ;
   U1015 : OAI22_X1 port map( A1 => n2153, A2 => n95, B1 => n2151, B2 => n92, 
                           ZN => n1005);
   U1016 : AOI221_X1 port map( B1 => n101, B2 => n3874, C1 => n98, C2 => n3908,
                           A => n1005, ZN => n1018);
   U1017 : OAI22_X1 port map( A1 => n2158, A2 => n107, B1 => n2156, B2 => n104,
                           ZN => n1008);
   U1018 : AOI221_X1 port map( B1 => n113, B2 => n4010, C1 => n110, C2 => n4044
                           , A => n1008, ZN => n1017);
   U1019 : OAI22_X1 port map( A1 => n2163, A2 => n119, B1 => n2161, B2 => n116,
                           ZN => n1011);
   U1020 : AOI221_X1 port map( B1 => n125, B2 => n4150, C1 => n122, C2 => n4185
                           , A => n1011, ZN => n1016);
   U1021 : OAI22_X1 port map( A1 => n2168, A2 => n131, B1 => n2166, B2 => n128,
                           ZN => n1014);
   U1022 : AOI221_X1 port map( B1 => n137, B2 => n4290, C1 => n134, C2 => n4356
                           , A => n1014, ZN => n1015);
   U1023 : NAND4_X1 port map( A1 => n1018, A2 => n1017, A3 => n1016, A4 => 
                           n1015, ZN => n1036);
   U1024 : OAI22_X1 port map( A1 => n2177, A2 => n143, B1 => n2175, B2 => n140,
                           ZN => n1021);
   U1025 : AOI221_X1 port map( B1 => n149, B2 => n2305, C1 => n146, C2 => n2339
                           , A => n1021, ZN => n1034);
   U1026 : OAI22_X1 port map( A1 => n2182, A2 => n155, B1 => n2180, B2 => n152,
                           ZN => n1024);
   U1027 : AOI221_X1 port map( B1 => n161, B2 => n2441, C1 => n158, C2 => n2479
                           , A => n1024, ZN => n1033);
   U1028 : OAI22_X1 port map( A1 => n2187, A2 => n167, B1 => n2185, B2 => n164,
                           ZN => n1027);
   U1029 : AOI221_X1 port map( B1 => n173, B2 => n2513, C1 => n170, C2 => n3635
                           , A => n1027, ZN => n1032);
   U1030 : OAI22_X1 port map( A1 => n2192, A2 => n179, B1 => n2190, B2 => n176,
                           ZN => n1030);
   U1031 : AOI221_X1 port map( B1 => n185, B2 => n3737, C1 => n182, C2 => n3771
                           , A => n1030, ZN => n1031);
   U1032 : NAND4_X1 port map( A1 => n1034, A2 => n1033, A3 => n1032, A4 => 
                           n1031, ZN => n1035);
   U1033 : OAI21_X1 port map( B1 => n1036, B2 => n1035, A => n188, ZN => n1037)
                           ;
   U1034 : OAI21_X1 port map( B1 => n191, B2 => n1038, A => n1037, ZN => n2558)
                           ;
   U1035 : OR2_X1 port map( A1 => RD1, A2 => n87, ZN => n2203);
   U1036 : INV_X1 port map( A => ADD_RD1(4), ZN => n1048);
   U1037 : INV_X1 port map( A => ADD_RD1(0), ZN => n1066);
   U1038 : INV_X1 port map( A => ADD_RD1(1), ZN => n1044);
   U1039 : NAND2_X1 port map( A1 => n74, A2 => n68, ZN => n2154);
   U1040 : NAND2_X1 port map( A1 => n75, A2 => n68, ZN => n2152);
   U1041 : OAI22_X1 port map( A1 => n195, A2 => n1041, B1 => n192, B2 => n1040,
                           ZN => n1042);
   U1042 : AOI221_X1 port map( B1 => n201, B2 => n3842, C1 => n198, C2 => n3876
                           , A => n1042, ZN => n1058);
   U1043 : INV_X1 port map( A => ADD_RD1(2), ZN => n1043);
   U1044 : NAND2_X1 port map( A1 => n74, A2 => n32, ZN => n2159);
   U1045 : NAND2_X1 port map( A1 => n75, A2 => n32, ZN => n2157);
   U1046 : OAI22_X1 port map( A1 => n207, A2 => n1046, B1 => n204, B2 => n1045,
                           ZN => n1047);
   U1047 : AOI221_X1 port map( B1 => n213, B2 => n3978, C1 => n210, C2 => n4012
                           , A => n1047, ZN => n1057);
   U1048 : INV_X1 port map( A => ADD_RD1(3), ZN => n1065);
   U1049 : NAND2_X1 port map( A1 => n73, A2 => n68, ZN => n2164);
   U1050 : NAND2_X1 port map( A1 => n35, A2 => n68, ZN => n2162);
   U1051 : OAI22_X1 port map( A1 => n219, A2 => n1050, B1 => n216, B2 => n1049,
                           ZN => n1051);
   U1052 : AOI221_X1 port map( B1 => n225, B2 => n4118, C1 => n222, C2 => n4153
                           , A => n1051, ZN => n1056);
   U1053 : NAND2_X1 port map( A1 => n73, A2 => n32, ZN => n2169);
   U1054 : NAND2_X1 port map( A1 => n35, A2 => n32, ZN => n2167);
   U1055 : OAI22_X1 port map( A1 => n231, A2 => n1053, B1 => n228, B2 => n1052,
                           ZN => n1054);
   U1056 : AOI221_X1 port map( B1 => n237, B2 => n4258, C1 => n234, C2 => n4293
                           , A => n1054, ZN => n1055);
   U1057 : NAND4_X1 port map( A1 => n1058, A2 => n1057, A3 => n1056, A4 => 
                           n1055, ZN => n1078);
   U1058 : NAND2_X1 port map( A1 => n3, A2 => n70, ZN => n2178);
   U1059 : NAND2_X1 port map( A1 => n3, A2 => n34, ZN => n2176);
   U1060 : OAI22_X1 port map( A1 => n243, A2 => n1060, B1 => n240, B2 => n1059,
                           ZN => n1061);
   U1061 : AOI221_X1 port map( B1 => n249, B2 => n2273, C1 => n246, C2 => n2307
                           , A => n1061, ZN => n1076);
   U1062 : NAND2_X1 port map( A1 => n4, A2 => n70, ZN => n2183);
   U1063 : NAND2_X1 port map( A1 => n4, A2 => n34, ZN => n2181);
   U1064 : OAI22_X1 port map( A1 => n255, A2 => n1063, B1 => n252, B2 => n1062,
                           ZN => n1064);
   U1065 : AOI221_X1 port map( B1 => n261, B2 => n2409, C1 => n258, C2 => n2447
                           , A => n1064, ZN => n1075);
   U1066 : NAND2_X1 port map( A1 => n80, A2 => n68, ZN => n2188);
   U1067 : NAND2_X1 port map( A1 => n79, A2 => n68, ZN => n2186);
   U1068 : OAI22_X1 port map( A1 => n267, A2 => n1068, B1 => n264, B2 => n1067,
                           ZN => n1069);
   U1069 : AOI221_X1 port map( B1 => n273, B2 => n2481, C1 => n270, C2 => n2515
                           , A => n1069, ZN => n1074);
   U1070 : NAND2_X1 port map( A1 => n80, A2 => n32, ZN => n2193);
   U1071 : NAND2_X1 port map( A1 => n79, A2 => n32, ZN => n2191);
   U1072 : OAI22_X1 port map( A1 => n279, A2 => n1071, B1 => n276, B2 => n1070,
                           ZN => n1072);
   U1073 : AOI221_X1 port map( B1 => n285, B2 => n3705, C1 => n282, C2 => n3739
                           , A => n1072, ZN => n1073);
   U1074 : NAND4_X1 port map( A1 => n1076, A2 => n1075, A3 => n1074, A4 => 
                           n1073, ZN => n1077);
   U1075 : OAI21_X1 port map( B1 => n1078, B2 => n1077, A => n288, ZN => n1079)
                           ;
   U1076 : OAI21_X1 port map( B1 => n291, B2 => n1080, A => n1079, ZN => n2559)
                           ;
   U1077 : OAI22_X1 port map( A1 => n195, A2 => n1082, B1 => n192, B2 => n1081,
                           ZN => n1083);
   U1078 : AOI221_X1 port map( B1 => n201, B2 => n3843, C1 => n198, C2 => n3877
                           , A => n1083, ZN => n1096);
   U1079 : OAI22_X1 port map( A1 => n207, A2 => n1085, B1 => n204, B2 => n1084,
                           ZN => n1086);
   U1080 : AOI221_X1 port map( B1 => n213, B2 => n3979, C1 => n210, C2 => n4013
                           , A => n1086, ZN => n1095);
   U1081 : OAI22_X1 port map( A1 => n219, A2 => n1088, B1 => n216, B2 => n1087,
                           ZN => n1089);
   U1082 : AOI221_X1 port map( B1 => n225, B2 => n4119, C1 => n222, C2 => n4154
                           , A => n1089, ZN => n1094);
   U1083 : OAI22_X1 port map( A1 => n231, A2 => n1091, B1 => n228, B2 => n1090,
                           ZN => n1092);
   U1084 : AOI221_X1 port map( B1 => n237, B2 => n4259, C1 => n234, C2 => n4295
                           , A => n1092, ZN => n1093);
   U1085 : NAND4_X1 port map( A1 => n1096, A2 => n1095, A3 => n1094, A4 => 
                           n1093, ZN => n1114);
   U1086 : OAI22_X1 port map( A1 => n243, A2 => n1098, B1 => n240, B2 => n1097,
                           ZN => n1099);
   U1087 : AOI221_X1 port map( B1 => n249, B2 => n2274, C1 => n246, C2 => n2308
                           , A => n1099, ZN => n1112);
   U1088 : OAI22_X1 port map( A1 => n255, A2 => n1101, B1 => n252, B2 => n1100,
                           ZN => n1102);
   U1089 : AOI221_X1 port map( B1 => n261, B2 => n2410, C1 => n258, C2 => n2448
                           , A => n1102, ZN => n1111);
   U1090 : OAI22_X1 port map( A1 => n267, A2 => n1104, B1 => n264, B2 => n1103,
                           ZN => n1105);
   U1091 : AOI221_X1 port map( B1 => n273, B2 => n2482, C1 => n270, C2 => n2516
                           , A => n1105, ZN => n1110);
   U1092 : OAI22_X1 port map( A1 => n279, A2 => n1107, B1 => n276, B2 => n1106,
                           ZN => n1108);
   U1093 : AOI221_X1 port map( B1 => n285, B2 => n3706, C1 => n282, C2 => n3740
                           , A => n1108, ZN => n1109);
   U1094 : NAND4_X1 port map( A1 => n1112, A2 => n1111, A3 => n1110, A4 => 
                           n1109, ZN => n1113);
   U1095 : OAI21_X1 port map( B1 => n1114, B2 => n1113, A => n288, ZN => n1115)
                           ;
   U1096 : OAI21_X1 port map( B1 => n291, B2 => n1116, A => n1115, ZN => n2560)
                           ;
   U1097 : OAI22_X1 port map( A1 => n195, A2 => n1118, B1 => n192, B2 => n1117,
                           ZN => n1119);
   U1098 : AOI221_X1 port map( B1 => n201, B2 => n3844, C1 => n198, C2 => n3878
                           , A => n1119, ZN => n1132);
   U1099 : OAI22_X1 port map( A1 => n207, A2 => n1121, B1 => n204, B2 => n1120,
                           ZN => n1122);
   U1100 : AOI221_X1 port map( B1 => n213, B2 => n3980, C1 => n210, C2 => n4014
                           , A => n1122, ZN => n1131);
   U1101 : OAI22_X1 port map( A1 => n219, A2 => n1124, B1 => n216, B2 => n1123,
                           ZN => n1125);
   U1102 : AOI221_X1 port map( B1 => n225, B2 => n4120, C1 => n222, C2 => n4155
                           , A => n1125, ZN => n1130);
   U1103 : OAI22_X1 port map( A1 => n231, A2 => n1127, B1 => n228, B2 => n1126,
                           ZN => n1128);
   U1104 : AOI221_X1 port map( B1 => n237, B2 => n4260, C1 => n234, C2 => n4297
                           , A => n1128, ZN => n1129);
   U1105 : NAND4_X1 port map( A1 => n1132, A2 => n1131, A3 => n1130, A4 => 
                           n1129, ZN => n1150);
   U1106 : OAI22_X1 port map( A1 => n243, A2 => n1134, B1 => n240, B2 => n1133,
                           ZN => n1135);
   U1107 : AOI221_X1 port map( B1 => n249, B2 => n2275, C1 => n246, C2 => n2309
                           , A => n1135, ZN => n1148);
   U1108 : OAI22_X1 port map( A1 => n255, A2 => n1137, B1 => n252, B2 => n1136,
                           ZN => n1138);
   U1109 : AOI221_X1 port map( B1 => n261, B2 => n2411, C1 => n258, C2 => n2449
                           , A => n1138, ZN => n1147);
   U1110 : OAI22_X1 port map( A1 => n267, A2 => n1140, B1 => n264, B2 => n1139,
                           ZN => n1141);
   U1111 : AOI221_X1 port map( B1 => n273, B2 => n2483, C1 => n270, C2 => n2517
                           , A => n1141, ZN => n1146);
   U1112 : OAI22_X1 port map( A1 => n279, A2 => n1143, B1 => n276, B2 => n1142,
                           ZN => n1144);
   U1113 : AOI221_X1 port map( B1 => n285, B2 => n3707, C1 => n282, C2 => n3741
                           , A => n1144, ZN => n1145);
   U1114 : NAND4_X1 port map( A1 => n1148, A2 => n1147, A3 => n1146, A4 => 
                           n1145, ZN => n1149);
   U1115 : OAI21_X1 port map( B1 => n1150, B2 => n1149, A => n288, ZN => n1151)
                           ;
   U1116 : OAI21_X1 port map( B1 => n291, B2 => n1152, A => n1151, ZN => n2561)
                           ;
   U1117 : OAI22_X1 port map( A1 => n195, A2 => n1154, B1 => n192, B2 => n1153,
                           ZN => n1155);
   U1118 : AOI221_X1 port map( B1 => n201, B2 => n3845, C1 => n198, C2 => n3879
                           , A => n1155, ZN => n1168);
   U1119 : OAI22_X1 port map( A1 => n207, A2 => n1157, B1 => n204, B2 => n1156,
                           ZN => n1158);
   U1120 : AOI221_X1 port map( B1 => n213, B2 => n3981, C1 => n210, C2 => n4015
                           , A => n1158, ZN => n1167);
   U1121 : OAI22_X1 port map( A1 => n219, A2 => n1160, B1 => n216, B2 => n1159,
                           ZN => n1161);
   U1122 : AOI221_X1 port map( B1 => n225, B2 => n4121, C1 => n222, C2 => n4156
                           , A => n1161, ZN => n1166);
   U1123 : OAI22_X1 port map( A1 => n231, A2 => n1163, B1 => n228, B2 => n1162,
                           ZN => n1164);
   U1124 : AOI221_X1 port map( B1 => n237, B2 => n4261, C1 => n234, C2 => n4299
                           , A => n1164, ZN => n1165);
   U1125 : NAND4_X1 port map( A1 => n1168, A2 => n1167, A3 => n1166, A4 => 
                           n1165, ZN => n1186);
   U1126 : OAI22_X1 port map( A1 => n243, A2 => n1170, B1 => n240, B2 => n1169,
                           ZN => n1171);
   U1127 : AOI221_X1 port map( B1 => n249, B2 => n2276, C1 => n246, C2 => n2310
                           , A => n1171, ZN => n1184);
   U1128 : OAI22_X1 port map( A1 => n255, A2 => n1173, B1 => n252, B2 => n1172,
                           ZN => n1174);
   U1129 : AOI221_X1 port map( B1 => n261, B2 => n2412, C1 => n258, C2 => n2450
                           , A => n1174, ZN => n1183);
   U1130 : OAI22_X1 port map( A1 => n267, A2 => n1176, B1 => n264, B2 => n1175,
                           ZN => n1177);
   U1131 : AOI221_X1 port map( B1 => n273, B2 => n2484, C1 => n270, C2 => n2518
                           , A => n1177, ZN => n1182);
   U1132 : OAI22_X1 port map( A1 => n279, A2 => n1179, B1 => n276, B2 => n1178,
                           ZN => n1180);
   U1133 : AOI221_X1 port map( B1 => n285, B2 => n3708, C1 => n282, C2 => n3742
                           , A => n1180, ZN => n1181);
   U1134 : NAND4_X1 port map( A1 => n1184, A2 => n1183, A3 => n1182, A4 => 
                           n1181, ZN => n1185);
   U1135 : OAI21_X1 port map( B1 => n1186, B2 => n1185, A => n288, ZN => n1187)
                           ;
   U1136 : OAI21_X1 port map( B1 => n291, B2 => n1188, A => n1187, ZN => n2562)
                           ;
   U1137 : OAI22_X1 port map( A1 => n195, A2 => n1190, B1 => n192, B2 => n1189,
                           ZN => n1191);
   U1138 : AOI221_X1 port map( B1 => n201, B2 => n3846, C1 => n198, C2 => n3880
                           , A => n1191, ZN => n1204);
   U1139 : OAI22_X1 port map( A1 => n207, A2 => n1193, B1 => n204, B2 => n1192,
                           ZN => n1194);
   U1140 : AOI221_X1 port map( B1 => n213, B2 => n3982, C1 => n210, C2 => n4016
                           , A => n1194, ZN => n1203);
   U1141 : OAI22_X1 port map( A1 => n219, A2 => n1196, B1 => n216, B2 => n1195,
                           ZN => n1197);
   U1142 : AOI221_X1 port map( B1 => n225, B2 => n4122, C1 => n222, C2 => n4157
                           , A => n1197, ZN => n1202);
   U1143 : OAI22_X1 port map( A1 => n231, A2 => n1199, B1 => n228, B2 => n1198,
                           ZN => n1200);
   U1144 : AOI221_X1 port map( B1 => n237, B2 => n4262, C1 => n234, C2 => n4301
                           , A => n1200, ZN => n1201);
   U1145 : NAND4_X1 port map( A1 => n1204, A2 => n1203, A3 => n1202, A4 => 
                           n1201, ZN => n1222);
   U1146 : OAI22_X1 port map( A1 => n243, A2 => n1206, B1 => n240, B2 => n1205,
                           ZN => n1207);
   U1147 : AOI221_X1 port map( B1 => n249, B2 => n2277, C1 => n246, C2 => n2311
                           , A => n1207, ZN => n1220);
   U1148 : OAI22_X1 port map( A1 => n255, A2 => n1209, B1 => n252, B2 => n1208,
                           ZN => n1210);
   U1149 : AOI221_X1 port map( B1 => n261, B2 => n2413, C1 => n258, C2 => n2451
                           , A => n1210, ZN => n1219);
   U1150 : OAI22_X1 port map( A1 => n267, A2 => n1212, B1 => n264, B2 => n1211,
                           ZN => n1213);
   U1151 : AOI221_X1 port map( B1 => n273, B2 => n2485, C1 => n270, C2 => n2519
                           , A => n1213, ZN => n1218);
   U1152 : OAI22_X1 port map( A1 => n279, A2 => n1215, B1 => n276, B2 => n1214,
                           ZN => n1216);
   U1153 : AOI221_X1 port map( B1 => n285, B2 => n3709, C1 => n282, C2 => n3743
                           , A => n1216, ZN => n1217);
   U1154 : NAND4_X1 port map( A1 => n1220, A2 => n1219, A3 => n1218, A4 => 
                           n1217, ZN => n1221);
   U1155 : OAI21_X1 port map( B1 => n1222, B2 => n1221, A => n288, ZN => n1223)
                           ;
   U1156 : OAI21_X1 port map( B1 => n291, B2 => n1224, A => n1223, ZN => n2563)
                           ;
   U1157 : OAI22_X1 port map( A1 => n195, A2 => n1226, B1 => n192, B2 => n1225,
                           ZN => n1227);
   U1158 : AOI221_X1 port map( B1 => n201, B2 => n3847, C1 => n198, C2 => n3881
                           , A => n1227, ZN => n1240);
   U1159 : OAI22_X1 port map( A1 => n207, A2 => n1229, B1 => n204, B2 => n1228,
                           ZN => n1230);
   U1160 : AOI221_X1 port map( B1 => n213, B2 => n3983, C1 => n210, C2 => n4017
                           , A => n1230, ZN => n1239);
   U1161 : OAI22_X1 port map( A1 => n219, A2 => n1232, B1 => n216, B2 => n1231,
                           ZN => n1233);
   U1162 : AOI221_X1 port map( B1 => n225, B2 => n4123, C1 => n222, C2 => n4158
                           , A => n1233, ZN => n1238);
   U1163 : OAI22_X1 port map( A1 => n231, A2 => n1235, B1 => n228, B2 => n1234,
                           ZN => n1236);
   U1164 : AOI221_X1 port map( B1 => n237, B2 => n4263, C1 => n234, C2 => n4303
                           , A => n1236, ZN => n1237);
   U1165 : NAND4_X1 port map( A1 => n1240, A2 => n1239, A3 => n1238, A4 => 
                           n1237, ZN => n1258);
   U1166 : OAI22_X1 port map( A1 => n243, A2 => n1242, B1 => n240, B2 => n1241,
                           ZN => n1243);
   U1167 : AOI221_X1 port map( B1 => n249, B2 => n2278, C1 => n246, C2 => n2312
                           , A => n1243, ZN => n1256);
   U1168 : OAI22_X1 port map( A1 => n255, A2 => n1245, B1 => n252, B2 => n1244,
                           ZN => n1246);
   U1169 : AOI221_X1 port map( B1 => n261, B2 => n2414, C1 => n258, C2 => n2452
                           , A => n1246, ZN => n1255);
   U1170 : OAI22_X1 port map( A1 => n267, A2 => n1248, B1 => n264, B2 => n1247,
                           ZN => n1249);
   U1171 : AOI221_X1 port map( B1 => n273, B2 => n2486, C1 => n270, C2 => n2520
                           , A => n1249, ZN => n1254);
   U1172 : OAI22_X1 port map( A1 => n279, A2 => n1251, B1 => n276, B2 => n1250,
                           ZN => n1252);
   U1173 : AOI221_X1 port map( B1 => n285, B2 => n3710, C1 => n282, C2 => n3744
                           , A => n1252, ZN => n1253);
   U1174 : NAND4_X1 port map( A1 => n1256, A2 => n1255, A3 => n1254, A4 => 
                           n1253, ZN => n1257);
   U1175 : OAI21_X1 port map( B1 => n1258, B2 => n1257, A => n288, ZN => n1259)
                           ;
   U1176 : OAI21_X1 port map( B1 => n291, B2 => n1260, A => n1259, ZN => n2564)
                           ;
   U1177 : OAI22_X1 port map( A1 => n195, A2 => n1262, B1 => n192, B2 => n1261,
                           ZN => n1263);
   U1178 : AOI221_X1 port map( B1 => n201, B2 => n3848, C1 => n198, C2 => n3882
                           , A => n1263, ZN => n1276);
   U1179 : OAI22_X1 port map( A1 => n207, A2 => n1265, B1 => n204, B2 => n1264,
                           ZN => n1266);
   U1180 : AOI221_X1 port map( B1 => n213, B2 => n3984, C1 => n210, C2 => n4018
                           , A => n1266, ZN => n1275);
   U1181 : OAI22_X1 port map( A1 => n219, A2 => n1268, B1 => n216, B2 => n1267,
                           ZN => n1269);
   U1182 : AOI221_X1 port map( B1 => n225, B2 => n4124, C1 => n222, C2 => n4159
                           , A => n1269, ZN => n1274);
   U1183 : OAI22_X1 port map( A1 => n231, A2 => n1271, B1 => n228, B2 => n1270,
                           ZN => n1272);
   U1184 : AOI221_X1 port map( B1 => n237, B2 => n4264, C1 => n234, C2 => n4305
                           , A => n1272, ZN => n1273);
   U1185 : NAND4_X1 port map( A1 => n1276, A2 => n1275, A3 => n1274, A4 => 
                           n1273, ZN => n1294);
   U1186 : OAI22_X1 port map( A1 => n243, A2 => n1278, B1 => n240, B2 => n1277,
                           ZN => n1279);
   U1187 : AOI221_X1 port map( B1 => n249, B2 => n2279, C1 => n246, C2 => n2313
                           , A => n1279, ZN => n1292);
   U1188 : OAI22_X1 port map( A1 => n255, A2 => n1281, B1 => n252, B2 => n1280,
                           ZN => n1282);
   U1189 : AOI221_X1 port map( B1 => n261, B2 => n2415, C1 => n258, C2 => n2453
                           , A => n1282, ZN => n1291);
   U1190 : OAI22_X1 port map( A1 => n267, A2 => n1284, B1 => n264, B2 => n1283,
                           ZN => n1285);
   U1191 : AOI221_X1 port map( B1 => n273, B2 => n2487, C1 => n270, C2 => n2521
                           , A => n1285, ZN => n1290);
   U1192 : OAI22_X1 port map( A1 => n279, A2 => n1287, B1 => n276, B2 => n1286,
                           ZN => n1288);
   U1193 : AOI221_X1 port map( B1 => n285, B2 => n3711, C1 => n282, C2 => n3745
                           , A => n1288, ZN => n1289);
   U1194 : NAND4_X1 port map( A1 => n1292, A2 => n1291, A3 => n1290, A4 => 
                           n1289, ZN => n1293);
   U1195 : OAI21_X1 port map( B1 => n1294, B2 => n1293, A => n288, ZN => n1295)
                           ;
   U1196 : OAI21_X1 port map( B1 => n291, B2 => n1296, A => n1295, ZN => n2565)
                           ;
   U1197 : OAI22_X1 port map( A1 => n195, A2 => n1298, B1 => n192, B2 => n1297,
                           ZN => n1299);
   U1198 : AOI221_X1 port map( B1 => n201, B2 => n3849, C1 => n198, C2 => n3883
                           , A => n1299, ZN => n1312);
   U1199 : OAI22_X1 port map( A1 => n207, A2 => n1301, B1 => n204, B2 => n1300,
                           ZN => n1302);
   U1200 : AOI221_X1 port map( B1 => n213, B2 => n3985, C1 => n210, C2 => n4019
                           , A => n1302, ZN => n1311);
   U1201 : OAI22_X1 port map( A1 => n219, A2 => n1304, B1 => n216, B2 => n1303,
                           ZN => n1305);
   U1202 : AOI221_X1 port map( B1 => n225, B2 => n4125, C1 => n222, C2 => n4160
                           , A => n1305, ZN => n1310);
   U1203 : OAI22_X1 port map( A1 => n231, A2 => n1307, B1 => n228, B2 => n1306,
                           ZN => n1308);
   U1204 : AOI221_X1 port map( B1 => n237, B2 => n4265, C1 => n234, C2 => n4307
                           , A => n1308, ZN => n1309);
   U1205 : NAND4_X1 port map( A1 => n1312, A2 => n1311, A3 => n1310, A4 => 
                           n1309, ZN => n1330);
   U1206 : OAI22_X1 port map( A1 => n243, A2 => n1314, B1 => n240, B2 => n1313,
                           ZN => n1315);
   U1207 : AOI221_X1 port map( B1 => n249, B2 => n2280, C1 => n246, C2 => n2314
                           , A => n1315, ZN => n1328);
   U1208 : OAI22_X1 port map( A1 => n255, A2 => n1317, B1 => n252, B2 => n1316,
                           ZN => n1318);
   U1209 : AOI221_X1 port map( B1 => n261, B2 => n2416, C1 => n258, C2 => n2454
                           , A => n1318, ZN => n1327);
   U1210 : OAI22_X1 port map( A1 => n267, A2 => n1320, B1 => n264, B2 => n1319,
                           ZN => n1321);
   U1211 : AOI221_X1 port map( B1 => n273, B2 => n2488, C1 => n270, C2 => n2522
                           , A => n1321, ZN => n1326);
   U1212 : OAI22_X1 port map( A1 => n279, A2 => n1323, B1 => n276, B2 => n1322,
                           ZN => n1324);
   U1213 : AOI221_X1 port map( B1 => n285, B2 => n3712, C1 => n282, C2 => n3746
                           , A => n1324, ZN => n1325);
   U1214 : NAND4_X1 port map( A1 => n1328, A2 => n1327, A3 => n1326, A4 => 
                           n1325, ZN => n1329);
   U1215 : OAI21_X1 port map( B1 => n1330, B2 => n1329, A => n288, ZN => n1331)
                           ;
   U1216 : OAI21_X1 port map( B1 => n291, B2 => n1332, A => n1331, ZN => n2566)
                           ;
   U1217 : OAI22_X1 port map( A1 => n195, A2 => n1334, B1 => n192, B2 => n1333,
                           ZN => n1335);
   U1218 : AOI221_X1 port map( B1 => n201, B2 => n3850, C1 => n198, C2 => n3884
                           , A => n1335, ZN => n1348);
   U1219 : OAI22_X1 port map( A1 => n207, A2 => n1337, B1 => n204, B2 => n1336,
                           ZN => n1338);
   U1220 : AOI221_X1 port map( B1 => n213, B2 => n3986, C1 => n210, C2 => n4020
                           , A => n1338, ZN => n1347);
   U1221 : OAI22_X1 port map( A1 => n219, A2 => n1340, B1 => n216, B2 => n1339,
                           ZN => n1341);
   U1222 : AOI221_X1 port map( B1 => n225, B2 => n4126, C1 => n222, C2 => n4161
                           , A => n1341, ZN => n1346);
   U1223 : OAI22_X1 port map( A1 => n231, A2 => n1343, B1 => n228, B2 => n1342,
                           ZN => n1344);
   U1224 : AOI221_X1 port map( B1 => n237, B2 => n4266, C1 => n234, C2 => n4309
                           , A => n1344, ZN => n1345);
   U1225 : NAND4_X1 port map( A1 => n1348, A2 => n1347, A3 => n1346, A4 => 
                           n1345, ZN => n1366);
   U1226 : OAI22_X1 port map( A1 => n243, A2 => n1350, B1 => n240, B2 => n1349,
                           ZN => n1351);
   U1227 : AOI221_X1 port map( B1 => n249, B2 => n2281, C1 => n246, C2 => n2315
                           , A => n1351, ZN => n1364);
   U1228 : OAI22_X1 port map( A1 => n255, A2 => n1353, B1 => n252, B2 => n1352,
                           ZN => n1354);
   U1229 : AOI221_X1 port map( B1 => n261, B2 => n2417, C1 => n258, C2 => n2455
                           , A => n1354, ZN => n1363);
   U1230 : OAI22_X1 port map( A1 => n267, A2 => n1356, B1 => n264, B2 => n1355,
                           ZN => n1357);
   U1231 : AOI221_X1 port map( B1 => n273, B2 => n2489, C1 => n270, C2 => n2523
                           , A => n1357, ZN => n1362);
   U1232 : OAI22_X1 port map( A1 => n279, A2 => n1359, B1 => n276, B2 => n1358,
                           ZN => n1360);
   U1233 : AOI221_X1 port map( B1 => n285, B2 => n3713, C1 => n282, C2 => n3747
                           , A => n1360, ZN => n1361);
   U1234 : NAND4_X1 port map( A1 => n1364, A2 => n1363, A3 => n1362, A4 => 
                           n1361, ZN => n1365);
   U1235 : OAI21_X1 port map( B1 => n1366, B2 => n1365, A => n288, ZN => n1367)
                           ;
   U1236 : OAI21_X1 port map( B1 => n291, B2 => n19, A => n1367, ZN => n2567);
   U1237 : OAI22_X1 port map( A1 => n195, A2 => n1369, B1 => n192, B2 => n1368,
                           ZN => n1370);
   U1238 : AOI221_X1 port map( B1 => n201, B2 => n3851, C1 => n198, C2 => n3885
                           , A => n1370, ZN => n1383);
   U1239 : OAI22_X1 port map( A1 => n207, A2 => n1372, B1 => n204, B2 => n1371,
                           ZN => n1373);
   U1240 : AOI221_X1 port map( B1 => n213, B2 => n3987, C1 => n210, C2 => n4021
                           , A => n1373, ZN => n1382);
   U1241 : OAI22_X1 port map( A1 => n219, A2 => n1375, B1 => n216, B2 => n1374,
                           ZN => n1376);
   U1242 : AOI221_X1 port map( B1 => n225, B2 => n4127, C1 => n222, C2 => n4162
                           , A => n1376, ZN => n1381);
   U1243 : OAI22_X1 port map( A1 => n231, A2 => n1378, B1 => n228, B2 => n1377,
                           ZN => n1379);
   U1244 : AOI221_X1 port map( B1 => n237, B2 => n4267, C1 => n234, C2 => n4311
                           , A => n1379, ZN => n1380);
   U1245 : NAND4_X1 port map( A1 => n1383, A2 => n1382, A3 => n1381, A4 => 
                           n1380, ZN => n1401);
   U1246 : OAI22_X1 port map( A1 => n243, A2 => n1385, B1 => n240, B2 => n1384,
                           ZN => n1386);
   U1247 : AOI221_X1 port map( B1 => n249, B2 => n2282, C1 => n246, C2 => n2316
                           , A => n1386, ZN => n1399);
   U1248 : OAI22_X1 port map( A1 => n255, A2 => n1388, B1 => n252, B2 => n1387,
                           ZN => n1389);
   U1249 : AOI221_X1 port map( B1 => n261, B2 => n2418, C1 => n258, C2 => n2456
                           , A => n1389, ZN => n1398);
   U1250 : OAI22_X1 port map( A1 => n267, A2 => n1391, B1 => n264, B2 => n1390,
                           ZN => n1392);
   U1251 : AOI221_X1 port map( B1 => n273, B2 => n2490, C1 => n270, C2 => n2524
                           , A => n1392, ZN => n1397);
   U1252 : OAI22_X1 port map( A1 => n279, A2 => n1394, B1 => n276, B2 => n1393,
                           ZN => n1395);
   U1253 : AOI221_X1 port map( B1 => n285, B2 => n3714, C1 => n282, C2 => n3748
                           , A => n1395, ZN => n1396);
   U1254 : NAND4_X1 port map( A1 => n1399, A2 => n1398, A3 => n1397, A4 => 
                           n1396, ZN => n1400);
   U1255 : OAI21_X1 port map( B1 => n1401, B2 => n1400, A => n288, ZN => n1402)
                           ;
   U1256 : OAI21_X1 port map( B1 => n291, B2 => n23, A => n1402, ZN => n2568);
   U1257 : OAI22_X1 port map( A1 => n195, A2 => n1404, B1 => n192, B2 => n1403,
                           ZN => n1405);
   U1258 : AOI221_X1 port map( B1 => n201, B2 => n3852, C1 => n198, C2 => n3886
                           , A => n1405, ZN => n1418);
   U1259 : OAI22_X1 port map( A1 => n207, A2 => n1407, B1 => n204, B2 => n1406,
                           ZN => n1408);
   U1260 : AOI221_X1 port map( B1 => n213, B2 => n3988, C1 => n210, C2 => n4022
                           , A => n1408, ZN => n1417);
   U1261 : OAI22_X1 port map( A1 => n219, A2 => n1410, B1 => n216, B2 => n1409,
                           ZN => n1411);
   U1262 : AOI221_X1 port map( B1 => n225, B2 => n4128, C1 => n222, C2 => n4163
                           , A => n1411, ZN => n1416);
   U1263 : OAI22_X1 port map( A1 => n231, A2 => n1413, B1 => n228, B2 => n1412,
                           ZN => n1414);
   U1264 : AOI221_X1 port map( B1 => n237, B2 => n4268, C1 => n234, C2 => n4313
                           , A => n1414, ZN => n1415);
   U1265 : NAND4_X1 port map( A1 => n1418, A2 => n1417, A3 => n1416, A4 => 
                           n1415, ZN => n1436);
   U1266 : OAI22_X1 port map( A1 => n243, A2 => n1420, B1 => n240, B2 => n1419,
                           ZN => n1421);
   U1267 : AOI221_X1 port map( B1 => n249, B2 => n2283, C1 => n246, C2 => n2317
                           , A => n1421, ZN => n1434);
   U1268 : OAI22_X1 port map( A1 => n255, A2 => n1423, B1 => n252, B2 => n1422,
                           ZN => n1424);
   U1269 : AOI221_X1 port map( B1 => n261, B2 => n2419, C1 => n258, C2 => n2457
                           , A => n1424, ZN => n1433);
   U1270 : OAI22_X1 port map( A1 => n267, A2 => n1426, B1 => n264, B2 => n1425,
                           ZN => n1427);
   U1271 : AOI221_X1 port map( B1 => n273, B2 => n2491, C1 => n270, C2 => n2525
                           , A => n1427, ZN => n1432);
   U1272 : OAI22_X1 port map( A1 => n279, A2 => n1429, B1 => n276, B2 => n1428,
                           ZN => n1430);
   U1273 : AOI221_X1 port map( B1 => n285, B2 => n3715, C1 => n282, C2 => n3749
                           , A => n1430, ZN => n1431);
   U1274 : NAND4_X1 port map( A1 => n1434, A2 => n1433, A3 => n1432, A4 => 
                           n1431, ZN => n1435);
   U1275 : OAI21_X1 port map( B1 => n1436, B2 => n1435, A => n288, ZN => n1437)
                           ;
   U1276 : OAI21_X1 port map( B1 => n291, B2 => n26, A => n1437, ZN => n2569);
   U1277 : OAI22_X1 port map( A1 => n195, A2 => n1439, B1 => n192, B2 => n1438,
                           ZN => n1440);
   U1278 : AOI221_X1 port map( B1 => n201, B2 => n3853, C1 => n198, C2 => n3887
                           , A => n1440, ZN => n1453);
   U1279 : OAI22_X1 port map( A1 => n207, A2 => n1442, B1 => n204, B2 => n1441,
                           ZN => n1443);
   U1280 : AOI221_X1 port map( B1 => n213, B2 => n3989, C1 => n210, C2 => n4023
                           , A => n1443, ZN => n1452);
   U1281 : OAI22_X1 port map( A1 => n219, A2 => n1445, B1 => n216, B2 => n1444,
                           ZN => n1446);
   U1282 : AOI221_X1 port map( B1 => n225, B2 => n4129, C1 => n222, C2 => n4164
                           , A => n1446, ZN => n1451);
   U1283 : OAI22_X1 port map( A1 => n231, A2 => n1448, B1 => n228, B2 => n1447,
                           ZN => n1449);
   U1284 : AOI221_X1 port map( B1 => n237, B2 => n4269, C1 => n234, C2 => n4315
                           , A => n1449, ZN => n1450);
   U1285 : NAND4_X1 port map( A1 => n1453, A2 => n1452, A3 => n1451, A4 => 
                           n1450, ZN => n1471);
   U1286 : OAI22_X1 port map( A1 => n243, A2 => n1455, B1 => n240, B2 => n1454,
                           ZN => n1456);
   U1287 : AOI221_X1 port map( B1 => n249, B2 => n2284, C1 => n246, C2 => n2318
                           , A => n1456, ZN => n1469);
   U1288 : OAI22_X1 port map( A1 => n255, A2 => n1458, B1 => n252, B2 => n1457,
                           ZN => n1459);
   U1289 : AOI221_X1 port map( B1 => n261, B2 => n2420, C1 => n258, C2 => n2458
                           , A => n1459, ZN => n1468);
   U1290 : OAI22_X1 port map( A1 => n267, A2 => n1461, B1 => n264, B2 => n1460,
                           ZN => n1462);
   U1291 : AOI221_X1 port map( B1 => n273, B2 => n2492, C1 => n270, C2 => n2526
                           , A => n1462, ZN => n1467);
   U1292 : OAI22_X1 port map( A1 => n279, A2 => n1464, B1 => n276, B2 => n1463,
                           ZN => n1465);
   U1293 : AOI221_X1 port map( B1 => n285, B2 => n3716, C1 => n282, C2 => n3750
                           , A => n1465, ZN => n1466);
   U1294 : NAND4_X1 port map( A1 => n1469, A2 => n1468, A3 => n1467, A4 => 
                           n1466, ZN => n1470);
   U1295 : OAI21_X1 port map( B1 => n1471, B2 => n1470, A => n288, ZN => n1472)
                           ;
   U1296 : OAI21_X1 port map( B1 => n292, B2 => n24, A => n1472, ZN => n2570);
   U1297 : OAI22_X1 port map( A1 => n196, A2 => n1474, B1 => n193, B2 => n1473,
                           ZN => n1475);
   U1298 : AOI221_X1 port map( B1 => n202, B2 => n3854, C1 => n199, C2 => n3888
                           , A => n1475, ZN => n1488);
   U1299 : OAI22_X1 port map( A1 => n208, A2 => n1477, B1 => n205, B2 => n1476,
                           ZN => n1478);
   U1300 : AOI221_X1 port map( B1 => n214, B2 => n3990, C1 => n211, C2 => n4024
                           , A => n1478, ZN => n1487);
   U1301 : OAI22_X1 port map( A1 => n220, A2 => n1480, B1 => n217, B2 => n1479,
                           ZN => n1481);
   U1302 : AOI221_X1 port map( B1 => n226, B2 => n4130, C1 => n223, C2 => n4165
                           , A => n1481, ZN => n1486);
   U1303 : OAI22_X1 port map( A1 => n232, A2 => n1483, B1 => n229, B2 => n1482,
                           ZN => n1484);
   U1304 : AOI221_X1 port map( B1 => n238, B2 => n4270, C1 => n235, C2 => n4317
                           , A => n1484, ZN => n1485);
   U1305 : NAND4_X1 port map( A1 => n1488, A2 => n1487, A3 => n1486, A4 => 
                           n1485, ZN => n1506);
   U1306 : OAI22_X1 port map( A1 => n244, A2 => n1490, B1 => n241, B2 => n1489,
                           ZN => n1491);
   U1307 : AOI221_X1 port map( B1 => n250, B2 => n2285, C1 => n247, C2 => n2319
                           , A => n1491, ZN => n1504);
   U1308 : OAI22_X1 port map( A1 => n256, A2 => n1493, B1 => n253, B2 => n1492,
                           ZN => n1494);
   U1309 : AOI221_X1 port map( B1 => n262, B2 => n2421, C1 => n259, C2 => n2459
                           , A => n1494, ZN => n1503);
   U1310 : OAI22_X1 port map( A1 => n268, A2 => n1496, B1 => n265, B2 => n1495,
                           ZN => n1497);
   U1311 : AOI221_X1 port map( B1 => n274, B2 => n2493, C1 => n271, C2 => n3615
                           , A => n1497, ZN => n1502);
   U1312 : OAI22_X1 port map( A1 => n280, A2 => n1499, B1 => n277, B2 => n1498,
                           ZN => n1500);
   U1313 : AOI221_X1 port map( B1 => n286, B2 => n3717, C1 => n283, C2 => n3751
                           , A => n1500, ZN => n1501);
   U1314 : NAND4_X1 port map( A1 => n1504, A2 => n1503, A3 => n1502, A4 => 
                           n1501, ZN => n1505);
   U1315 : OAI21_X1 port map( B1 => n1506, B2 => n1505, A => n289, ZN => n1507)
                           ;
   U1316 : OAI21_X1 port map( B1 => n292, B2 => n25, A => n1507, ZN => n2571);
   U1317 : OAI22_X1 port map( A1 => n196, A2 => n1509, B1 => n193, B2 => n1508,
                           ZN => n1510);
   U1318 : AOI221_X1 port map( B1 => n202, B2 => n3855, C1 => n199, C2 => n3889
                           , A => n1510, ZN => n1523);
   U1319 : OAI22_X1 port map( A1 => n208, A2 => n1512, B1 => n205, B2 => n1511,
                           ZN => n1513);
   U1320 : AOI221_X1 port map( B1 => n214, B2 => n3991, C1 => n211, C2 => n4025
                           , A => n1513, ZN => n1522);
   U1321 : OAI22_X1 port map( A1 => n220, A2 => n1515, B1 => n217, B2 => n1514,
                           ZN => n1516);
   U1322 : AOI221_X1 port map( B1 => n226, B2 => n4131, C1 => n223, C2 => n4166
                           , A => n1516, ZN => n1521);
   U1323 : OAI22_X1 port map( A1 => n232, A2 => n1518, B1 => n229, B2 => n1517,
                           ZN => n1519);
   U1324 : AOI221_X1 port map( B1 => n238, B2 => n4271, C1 => n235, C2 => n4319
                           , A => n1519, ZN => n1520);
   U1325 : NAND4_X1 port map( A1 => n1523, A2 => n1522, A3 => n1521, A4 => 
                           n1520, ZN => n1541);
   U1326 : OAI22_X1 port map( A1 => n244, A2 => n1525, B1 => n241, B2 => n1524,
                           ZN => n1526);
   U1327 : AOI221_X1 port map( B1 => n250, B2 => n2286, C1 => n247, C2 => n2320
                           , A => n1526, ZN => n1539);
   U1328 : OAI22_X1 port map( A1 => n256, A2 => n1528, B1 => n253, B2 => n1527,
                           ZN => n1529);
   U1329 : AOI221_X1 port map( B1 => n262, B2 => n2422, C1 => n259, C2 => n2460
                           , A => n1529, ZN => n1538);
   U1330 : OAI22_X1 port map( A1 => n268, A2 => n1531, B1 => n265, B2 => n1530,
                           ZN => n1532);
   U1331 : AOI221_X1 port map( B1 => n274, B2 => n2494, C1 => n271, C2 => n3616
                           , A => n1532, ZN => n1537);
   U1332 : OAI22_X1 port map( A1 => n280, A2 => n1534, B1 => n277, B2 => n1533,
                           ZN => n1535);
   U1333 : AOI221_X1 port map( B1 => n286, B2 => n3718, C1 => n283, C2 => n3752
                           , A => n1535, ZN => n1536);
   U1334 : NAND4_X1 port map( A1 => n1539, A2 => n1538, A3 => n1537, A4 => 
                           n1536, ZN => n1540);
   U1335 : OAI21_X1 port map( B1 => n1541, B2 => n1540, A => n289, ZN => n1542)
                           ;
   U1336 : OAI21_X1 port map( B1 => n292, B2 => n1543, A => n1542, ZN => n2572)
                           ;
   U1337 : OAI22_X1 port map( A1 => n196, A2 => n1545, B1 => n193, B2 => n1544,
                           ZN => n1546);
   U1338 : AOI221_X1 port map( B1 => n202, B2 => n3856, C1 => n199, C2 => n3890
                           , A => n1546, ZN => n1559);
   U1339 : OAI22_X1 port map( A1 => n208, A2 => n1548, B1 => n205, B2 => n1547,
                           ZN => n1549);
   U1340 : AOI221_X1 port map( B1 => n214, B2 => n3992, C1 => n211, C2 => n4026
                           , A => n1549, ZN => n1558);
   U1341 : OAI22_X1 port map( A1 => n220, A2 => n1551, B1 => n217, B2 => n1550,
                           ZN => n1552);
   U1342 : AOI221_X1 port map( B1 => n226, B2 => n4132, C1 => n223, C2 => n4167
                           , A => n1552, ZN => n1557);
   U1343 : OAI22_X1 port map( A1 => n232, A2 => n1554, B1 => n229, B2 => n1553,
                           ZN => n1555);
   U1344 : AOI221_X1 port map( B1 => n238, B2 => n4272, C1 => n235, C2 => n4321
                           , A => n1555, ZN => n1556);
   U1345 : NAND4_X1 port map( A1 => n1559, A2 => n1558, A3 => n1557, A4 => 
                           n1556, ZN => n1577);
   U1346 : OAI22_X1 port map( A1 => n244, A2 => n1561, B1 => n241, B2 => n1560,
                           ZN => n1562);
   U1347 : AOI221_X1 port map( B1 => n250, B2 => n2287, C1 => n247, C2 => n2321
                           , A => n1562, ZN => n1575);
   U1348 : OAI22_X1 port map( A1 => n256, A2 => n1564, B1 => n253, B2 => n1563,
                           ZN => n1565);
   U1349 : AOI221_X1 port map( B1 => n262, B2 => n2423, C1 => n259, C2 => n2461
                           , A => n1565, ZN => n1574);
   U1350 : OAI22_X1 port map( A1 => n268, A2 => n1567, B1 => n265, B2 => n1566,
                           ZN => n1568);
   U1351 : AOI221_X1 port map( B1 => n274, B2 => n2495, C1 => n271, C2 => n3617
                           , A => n1568, ZN => n1573);
   U1352 : OAI22_X1 port map( A1 => n280, A2 => n1570, B1 => n277, B2 => n1569,
                           ZN => n1571);
   U1353 : AOI221_X1 port map( B1 => n286, B2 => n3719, C1 => n283, C2 => n3753
                           , A => n1571, ZN => n1572);
   U1354 : NAND4_X1 port map( A1 => n1575, A2 => n1574, A3 => n1573, A4 => 
                           n1572, ZN => n1576);
   U1355 : OAI21_X1 port map( B1 => n1577, B2 => n1576, A => n289, ZN => n1578)
                           ;
   U1356 : OAI21_X1 port map( B1 => n292, B2 => n21, A => n1578, ZN => n2573);
   U1357 : OAI22_X1 port map( A1 => n196, A2 => n1580, B1 => n193, B2 => n1579,
                           ZN => n1581);
   U1358 : AOI221_X1 port map( B1 => n202, B2 => n3857, C1 => n199, C2 => n3891
                           , A => n1581, ZN => n1594);
   U1359 : OAI22_X1 port map( A1 => n208, A2 => n1583, B1 => n205, B2 => n1582,
                           ZN => n1584);
   U1360 : AOI221_X1 port map( B1 => n214, B2 => n3993, C1 => n211, C2 => n4027
                           , A => n1584, ZN => n1593);
   U1361 : OAI22_X1 port map( A1 => n220, A2 => n1586, B1 => n217, B2 => n1585,
                           ZN => n1587);
   U1362 : AOI221_X1 port map( B1 => n226, B2 => n4133, C1 => n223, C2 => n4168
                           , A => n1587, ZN => n1592);
   U1363 : OAI22_X1 port map( A1 => n232, A2 => n1589, B1 => n229, B2 => n1588,
                           ZN => n1590);
   U1364 : AOI221_X1 port map( B1 => n238, B2 => n4273, C1 => n235, C2 => n4323
                           , A => n1590, ZN => n1591);
   U1365 : NAND4_X1 port map( A1 => n1594, A2 => n1593, A3 => n1592, A4 => 
                           n1591, ZN => n1612);
   U1366 : OAI22_X1 port map( A1 => n244, A2 => n1596, B1 => n241, B2 => n1595,
                           ZN => n1597);
   U1367 : AOI221_X1 port map( B1 => n250, B2 => n2288, C1 => n247, C2 => n2322
                           , A => n1597, ZN => n1610);
   U1368 : OAI22_X1 port map( A1 => n256, A2 => n1599, B1 => n253, B2 => n1598,
                           ZN => n1600);
   U1369 : AOI221_X1 port map( B1 => n262, B2 => n2424, C1 => n259, C2 => n2462
                           , A => n1600, ZN => n1609);
   U1370 : OAI22_X1 port map( A1 => n268, A2 => n1602, B1 => n265, B2 => n1601,
                           ZN => n1603);
   U1371 : AOI221_X1 port map( B1 => n274, B2 => n2496, C1 => n271, C2 => n3618
                           , A => n1603, ZN => n1608);
   U1372 : OAI22_X1 port map( A1 => n280, A2 => n1605, B1 => n277, B2 => n1604,
                           ZN => n1606);
   U1373 : AOI221_X1 port map( B1 => n286, B2 => n3720, C1 => n283, C2 => n3754
                           , A => n1606, ZN => n1607);
   U1374 : NAND4_X1 port map( A1 => n1610, A2 => n1609, A3 => n1608, A4 => 
                           n1607, ZN => n1611);
   U1375 : OAI21_X1 port map( B1 => n1612, B2 => n1611, A => n289, ZN => n1613)
                           ;
   U1376 : OAI21_X1 port map( B1 => n292, B2 => n22, A => n1613, ZN => n2574);
   U1377 : OAI22_X1 port map( A1 => n196, A2 => n1615, B1 => n193, B2 => n1614,
                           ZN => n1616);
   U1378 : AOI221_X1 port map( B1 => n202, B2 => n3858, C1 => n199, C2 => n3892
                           , A => n1616, ZN => n1629);
   U1379 : OAI22_X1 port map( A1 => n208, A2 => n1618, B1 => n205, B2 => n1617,
                           ZN => n1619);
   U1380 : AOI221_X1 port map( B1 => n214, B2 => n3994, C1 => n211, C2 => n4028
                           , A => n1619, ZN => n1628);
   U1381 : OAI22_X1 port map( A1 => n220, A2 => n1621, B1 => n217, B2 => n1620,
                           ZN => n1622);
   U1382 : AOI221_X1 port map( B1 => n226, B2 => n4134, C1 => n223, C2 => n4169
                           , A => n1622, ZN => n1627);
   U1383 : OAI22_X1 port map( A1 => n232, A2 => n1624, B1 => n229, B2 => n1623,
                           ZN => n1625);
   U1384 : AOI221_X1 port map( B1 => n238, B2 => n4274, C1 => n235, C2 => n4325
                           , A => n1625, ZN => n1626);
   U1385 : NAND4_X1 port map( A1 => n1629, A2 => n1628, A3 => n1627, A4 => 
                           n1626, ZN => n1647);
   U1386 : OAI22_X1 port map( A1 => n244, A2 => n1631, B1 => n241, B2 => n1630,
                           ZN => n1632);
   U1387 : AOI221_X1 port map( B1 => n250, B2 => n2289, C1 => n247, C2 => n2323
                           , A => n1632, ZN => n1645);
   U1388 : OAI22_X1 port map( A1 => n256, A2 => n1634, B1 => n253, B2 => n1633,
                           ZN => n1635);
   U1389 : AOI221_X1 port map( B1 => n262, B2 => n2425, C1 => n259, C2 => n2463
                           , A => n1635, ZN => n1644);
   U1390 : OAI22_X1 port map( A1 => n268, A2 => n1637, B1 => n265, B2 => n1636,
                           ZN => n1638);
   U1391 : AOI221_X1 port map( B1 => n274, B2 => n2497, C1 => n271, C2 => n3619
                           , A => n1638, ZN => n1643);
   U1392 : OAI22_X1 port map( A1 => n280, A2 => n1640, B1 => n277, B2 => n1639,
                           ZN => n1641);
   U1393 : AOI221_X1 port map( B1 => n286, B2 => n3721, C1 => n283, C2 => n3755
                           , A => n1641, ZN => n1642);
   U1394 : NAND4_X1 port map( A1 => n1645, A2 => n1644, A3 => n1643, A4 => 
                           n1642, ZN => n1646);
   U1395 : OAI21_X1 port map( B1 => n1647, B2 => n1646, A => n289, ZN => n1648)
                           ;
   U1396 : OAI21_X1 port map( B1 => n292, B2 => n1649, A => n1648, ZN => n2575)
                           ;
   U1397 : OAI22_X1 port map( A1 => n196, A2 => n1651, B1 => n193, B2 => n1650,
                           ZN => n1652);
   U1398 : AOI221_X1 port map( B1 => n202, B2 => n3859, C1 => n199, C2 => n3893
                           , A => n1652, ZN => n1665);
   U1399 : OAI22_X1 port map( A1 => n208, A2 => n1654, B1 => n205, B2 => n1653,
                           ZN => n1655);
   U1400 : AOI221_X1 port map( B1 => n214, B2 => n3995, C1 => n211, C2 => n4029
                           , A => n1655, ZN => n1664);
   U1401 : OAI22_X1 port map( A1 => n220, A2 => n1657, B1 => n217, B2 => n1656,
                           ZN => n1658);
   U1402 : AOI221_X1 port map( B1 => n226, B2 => n4135, C1 => n223, C2 => n4170
                           , A => n1658, ZN => n1663);
   U1403 : OAI22_X1 port map( A1 => n232, A2 => n1660, B1 => n229, B2 => n1659,
                           ZN => n1661);
   U1404 : AOI221_X1 port map( B1 => n238, B2 => n4275, C1 => n235, C2 => n4327
                           , A => n1661, ZN => n1662);
   U1405 : NAND4_X1 port map( A1 => n1665, A2 => n1664, A3 => n1663, A4 => 
                           n1662, ZN => n1683);
   U1406 : OAI22_X1 port map( A1 => n244, A2 => n1667, B1 => n241, B2 => n1666,
                           ZN => n1668);
   U1407 : AOI221_X1 port map( B1 => n250, B2 => n2290, C1 => n247, C2 => n2324
                           , A => n1668, ZN => n1681);
   U1408 : OAI22_X1 port map( A1 => n256, A2 => n1670, B1 => n253, B2 => n1669,
                           ZN => n1671);
   U1409 : AOI221_X1 port map( B1 => n262, B2 => n2426, C1 => n259, C2 => n2464
                           , A => n1671, ZN => n1680);
   U1410 : OAI22_X1 port map( A1 => n268, A2 => n1673, B1 => n265, B2 => n1672,
                           ZN => n1674);
   U1411 : AOI221_X1 port map( B1 => n274, B2 => n2498, C1 => n271, C2 => n3620
                           , A => n1674, ZN => n1679);
   U1412 : OAI22_X1 port map( A1 => n280, A2 => n1676, B1 => n277, B2 => n1675,
                           ZN => n1677);
   U1413 : AOI221_X1 port map( B1 => n286, B2 => n3722, C1 => n283, C2 => n3756
                           , A => n1677, ZN => n1678);
   U1414 : NAND4_X1 port map( A1 => n1681, A2 => n1680, A3 => n1679, A4 => 
                           n1678, ZN => n1682);
   U1415 : OAI21_X1 port map( B1 => n1683, B2 => n1682, A => n289, ZN => n1684)
                           ;
   U1416 : OAI21_X1 port map( B1 => n292, B2 => n1685, A => n1684, ZN => n2576)
                           ;
   U1417 : OAI22_X1 port map( A1 => n196, A2 => n1687, B1 => n193, B2 => n1686,
                           ZN => n1688);
   U1418 : AOI221_X1 port map( B1 => n202, B2 => n3860, C1 => n199, C2 => n3894
                           , A => n1688, ZN => n1701);
   U1419 : OAI22_X1 port map( A1 => n208, A2 => n1690, B1 => n205, B2 => n1689,
                           ZN => n1691);
   U1420 : AOI221_X1 port map( B1 => n214, B2 => n3996, C1 => n211, C2 => n4030
                           , A => n1691, ZN => n1700);
   U1421 : OAI22_X1 port map( A1 => n220, A2 => n1693, B1 => n217, B2 => n1692,
                           ZN => n1694);
   U1422 : AOI221_X1 port map( B1 => n226, B2 => n4136, C1 => n223, C2 => n4171
                           , A => n1694, ZN => n1699);
   U1423 : OAI22_X1 port map( A1 => n232, A2 => n1696, B1 => n229, B2 => n1695,
                           ZN => n1697);
   U1424 : AOI221_X1 port map( B1 => n238, B2 => n4276, C1 => n235, C2 => n4329
                           , A => n1697, ZN => n1698);
   U1425 : NAND4_X1 port map( A1 => n1701, A2 => n1700, A3 => n1699, A4 => 
                           n1698, ZN => n1719);
   U1426 : OAI22_X1 port map( A1 => n244, A2 => n1703, B1 => n241, B2 => n1702,
                           ZN => n1704);
   U1427 : AOI221_X1 port map( B1 => n250, B2 => n2291, C1 => n247, C2 => n2325
                           , A => n1704, ZN => n1717);
   U1428 : OAI22_X1 port map( A1 => n256, A2 => n1706, B1 => n253, B2 => n1705,
                           ZN => n1707);
   U1429 : AOI221_X1 port map( B1 => n262, B2 => n2427, C1 => n259, C2 => n2465
                           , A => n1707, ZN => n1716);
   U1430 : OAI22_X1 port map( A1 => n268, A2 => n1709, B1 => n265, B2 => n1708,
                           ZN => n1710);
   U1431 : AOI221_X1 port map( B1 => n274, B2 => n2499, C1 => n271, C2 => n3621
                           , A => n1710, ZN => n1715);
   U1432 : OAI22_X1 port map( A1 => n280, A2 => n1712, B1 => n277, B2 => n1711,
                           ZN => n1713);
   U1433 : AOI221_X1 port map( B1 => n286, B2 => n3723, C1 => n283, C2 => n3757
                           , A => n1713, ZN => n1714);
   U1434 : NAND4_X1 port map( A1 => n1717, A2 => n1716, A3 => n1715, A4 => 
                           n1714, ZN => n1718);
   U1435 : OAI21_X1 port map( B1 => n1719, B2 => n1718, A => n289, ZN => n1720)
                           ;
   U1436 : OAI21_X1 port map( B1 => n292, B2 => n17, A => n1720, ZN => n2577);
   U1437 : OAI22_X1 port map( A1 => n196, A2 => n1722, B1 => n193, B2 => n1721,
                           ZN => n1723);
   U1438 : AOI221_X1 port map( B1 => n202, B2 => n3861, C1 => n199, C2 => n3895
                           , A => n1723, ZN => n1736);
   U1439 : OAI22_X1 port map( A1 => n208, A2 => n1725, B1 => n205, B2 => n1724,
                           ZN => n1726);
   U1440 : AOI221_X1 port map( B1 => n214, B2 => n3997, C1 => n211, C2 => n4031
                           , A => n1726, ZN => n1735);
   U1441 : OAI22_X1 port map( A1 => n220, A2 => n1728, B1 => n217, B2 => n1727,
                           ZN => n1729);
   U1442 : AOI221_X1 port map( B1 => n226, B2 => n4137, C1 => n223, C2 => n4172
                           , A => n1729, ZN => n1734);
   U1443 : OAI22_X1 port map( A1 => n232, A2 => n1731, B1 => n229, B2 => n1730,
                           ZN => n1732);
   U1444 : AOI221_X1 port map( B1 => n238, B2 => n4277, C1 => n235, C2 => n4331
                           , A => n1732, ZN => n1733);
   U1445 : NAND4_X1 port map( A1 => n1736, A2 => n1735, A3 => n1734, A4 => 
                           n1733, ZN => n1754);
   U1446 : OAI22_X1 port map( A1 => n244, A2 => n1738, B1 => n241, B2 => n1737,
                           ZN => n1739);
   U1447 : AOI221_X1 port map( B1 => n250, B2 => n2292, C1 => n247, C2 => n2326
                           , A => n1739, ZN => n1752);
   U1448 : OAI22_X1 port map( A1 => n256, A2 => n1741, B1 => n253, B2 => n1740,
                           ZN => n1742);
   U1449 : AOI221_X1 port map( B1 => n262, B2 => n2428, C1 => n259, C2 => n2466
                           , A => n1742, ZN => n1751);
   U1450 : OAI22_X1 port map( A1 => n268, A2 => n1744, B1 => n265, B2 => n1743,
                           ZN => n1745);
   U1451 : AOI221_X1 port map( B1 => n274, B2 => n2500, C1 => n271, C2 => n3622
                           , A => n1745, ZN => n1750);
   U1452 : OAI22_X1 port map( A1 => n280, A2 => n1747, B1 => n277, B2 => n1746,
                           ZN => n1748);
   U1453 : AOI221_X1 port map( B1 => n286, B2 => n3724, C1 => n283, C2 => n3758
                           , A => n1748, ZN => n1749);
   U1454 : NAND4_X1 port map( A1 => n1752, A2 => n1751, A3 => n1750, A4 => 
                           n1749, ZN => n1753);
   U1455 : OAI21_X1 port map( B1 => n1754, B2 => n1753, A => n289, ZN => n1755)
                           ;
   U1456 : OAI21_X1 port map( B1 => n292, B2 => n1756, A => n1755, ZN => n2578)
                           ;
   U1457 : OAI22_X1 port map( A1 => n196, A2 => n1758, B1 => n193, B2 => n1757,
                           ZN => n1759);
   U1458 : AOI221_X1 port map( B1 => n202, B2 => n3862, C1 => n199, C2 => n3896
                           , A => n1759, ZN => n1772);
   U1459 : OAI22_X1 port map( A1 => n208, A2 => n1761, B1 => n205, B2 => n1760,
                           ZN => n1762);
   U1460 : AOI221_X1 port map( B1 => n214, B2 => n3998, C1 => n211, C2 => n4032
                           , A => n1762, ZN => n1771);
   U1461 : OAI22_X1 port map( A1 => n220, A2 => n1764, B1 => n217, B2 => n1763,
                           ZN => n1765);
   U1462 : AOI221_X1 port map( B1 => n226, B2 => n4138, C1 => n223, C2 => n4173
                           , A => n1765, ZN => n1770);
   U1463 : OAI22_X1 port map( A1 => n232, A2 => n1767, B1 => n229, B2 => n1766,
                           ZN => n1768);
   U1464 : AOI221_X1 port map( B1 => n238, B2 => n4278, C1 => n235, C2 => n4333
                           , A => n1768, ZN => n1769);
   U1465 : NAND4_X1 port map( A1 => n1772, A2 => n1771, A3 => n1770, A4 => 
                           n1769, ZN => n1790);
   U1466 : OAI22_X1 port map( A1 => n244, A2 => n1774, B1 => n241, B2 => n1773,
                           ZN => n1775);
   U1467 : AOI221_X1 port map( B1 => n250, B2 => n2293, C1 => n247, C2 => n2327
                           , A => n1775, ZN => n1788);
   U1468 : OAI22_X1 port map( A1 => n256, A2 => n1777, B1 => n253, B2 => n1776,
                           ZN => n1778);
   U1469 : AOI221_X1 port map( B1 => n262, B2 => n2429, C1 => n259, C2 => n2467
                           , A => n1778, ZN => n1787);
   U1470 : OAI22_X1 port map( A1 => n268, A2 => n1780, B1 => n265, B2 => n1779,
                           ZN => n1781);
   U1471 : AOI221_X1 port map( B1 => n274, B2 => n2501, C1 => n271, C2 => n3623
                           , A => n1781, ZN => n1786);
   U1472 : OAI22_X1 port map( A1 => n280, A2 => n1783, B1 => n277, B2 => n1782,
                           ZN => n1784);
   U1473 : AOI221_X1 port map( B1 => n286, B2 => n3725, C1 => n283, C2 => n3759
                           , A => n1784, ZN => n1785);
   U1474 : NAND4_X1 port map( A1 => n1788, A2 => n1787, A3 => n1786, A4 => 
                           n1785, ZN => n1789);
   U1475 : OAI21_X1 port map( B1 => n1790, B2 => n1789, A => n289, ZN => n1791)
                           ;
   U1476 : OAI21_X1 port map( B1 => n292, B2 => n1792, A => n1791, ZN => n2579)
                           ;
   U1477 : OAI22_X1 port map( A1 => n196, A2 => n1794, B1 => n193, B2 => n1793,
                           ZN => n1795);
   U1478 : AOI221_X1 port map( B1 => n202, B2 => n3863, C1 => n199, C2 => n3897
                           , A => n1795, ZN => n1808);
   U1479 : OAI22_X1 port map( A1 => n208, A2 => n1797, B1 => n205, B2 => n1796,
                           ZN => n1798);
   U1480 : AOI221_X1 port map( B1 => n214, B2 => n3999, C1 => n211, C2 => n4033
                           , A => n1798, ZN => n1807);
   U1481 : OAI22_X1 port map( A1 => n220, A2 => n1800, B1 => n217, B2 => n1799,
                           ZN => n1801);
   U1482 : AOI221_X1 port map( B1 => n226, B2 => n4139, C1 => n223, C2 => n4174
                           , A => n1801, ZN => n1806);
   U1483 : OAI22_X1 port map( A1 => n232, A2 => n1803, B1 => n229, B2 => n1802,
                           ZN => n1804);
   U1484 : AOI221_X1 port map( B1 => n238, B2 => n4279, C1 => n235, C2 => n4335
                           , A => n1804, ZN => n1805);
   U1485 : NAND4_X1 port map( A1 => n1808, A2 => n1807, A3 => n1806, A4 => 
                           n1805, ZN => n1826);
   U1486 : OAI22_X1 port map( A1 => n244, A2 => n1810, B1 => n241, B2 => n1809,
                           ZN => n1811);
   U1487 : AOI221_X1 port map( B1 => n250, B2 => n2294, C1 => n247, C2 => n2328
                           , A => n1811, ZN => n1824);
   U1488 : OAI22_X1 port map( A1 => n256, A2 => n1813, B1 => n253, B2 => n1812,
                           ZN => n1814);
   U1489 : AOI221_X1 port map( B1 => n262, B2 => n2430, C1 => n259, C2 => n2468
                           , A => n1814, ZN => n1823);
   U1490 : OAI22_X1 port map( A1 => n268, A2 => n1816, B1 => n265, B2 => n1815,
                           ZN => n1817);
   U1491 : AOI221_X1 port map( B1 => n274, B2 => n2502, C1 => n271, C2 => n3624
                           , A => n1817, ZN => n1822);
   U1492 : OAI22_X1 port map( A1 => n280, A2 => n1819, B1 => n277, B2 => n1818,
                           ZN => n1820);
   U1493 : AOI221_X1 port map( B1 => n286, B2 => n3726, C1 => n283, C2 => n3760
                           , A => n1820, ZN => n1821);
   U1494 : NAND4_X1 port map( A1 => n1824, A2 => n1823, A3 => n1822, A4 => 
                           n1821, ZN => n1825);
   U1495 : OAI21_X1 port map( B1 => n1826, B2 => n1825, A => n289, ZN => n1827)
                           ;
   U1496 : OAI21_X1 port map( B1 => n292, B2 => n1828, A => n1827, ZN => n2580)
                           ;
   U1497 : OAI22_X1 port map( A1 => n196, A2 => n1830, B1 => n193, B2 => n1829,
                           ZN => n1831);
   U1498 : AOI221_X1 port map( B1 => n202, B2 => n3864, C1 => n199, C2 => n3898
                           , A => n1831, ZN => n1844);
   U1499 : OAI22_X1 port map( A1 => n208, A2 => n1833, B1 => n205, B2 => n1832,
                           ZN => n1834);
   U1500 : AOI221_X1 port map( B1 => n214, B2 => n4000, C1 => n211, C2 => n4034
                           , A => n1834, ZN => n1843);
   U1501 : OAI22_X1 port map( A1 => n220, A2 => n1836, B1 => n217, B2 => n1835,
                           ZN => n1837);
   U1502 : AOI221_X1 port map( B1 => n226, B2 => n4140, C1 => n223, C2 => n4175
                           , A => n1837, ZN => n1842);
   U1503 : OAI22_X1 port map( A1 => n232, A2 => n1839, B1 => n229, B2 => n1838,
                           ZN => n1840);
   U1504 : AOI221_X1 port map( B1 => n238, B2 => n4280, C1 => n235, C2 => n4337
                           , A => n1840, ZN => n1841);
   U1505 : NAND4_X1 port map( A1 => n1844, A2 => n1843, A3 => n1842, A4 => 
                           n1841, ZN => n1862);
   U1506 : OAI22_X1 port map( A1 => n244, A2 => n1846, B1 => n241, B2 => n1845,
                           ZN => n1847);
   U1507 : AOI221_X1 port map( B1 => n250, B2 => n2295, C1 => n247, C2 => n2329
                           , A => n1847, ZN => n1860);
   U1508 : OAI22_X1 port map( A1 => n256, A2 => n1849, B1 => n253, B2 => n1848,
                           ZN => n1850);
   U1509 : AOI221_X1 port map( B1 => n262, B2 => n2431, C1 => n259, C2 => n2469
                           , A => n1850, ZN => n1859);
   U1510 : OAI22_X1 port map( A1 => n268, A2 => n1852, B1 => n265, B2 => n1851,
                           ZN => n1853);
   U1511 : AOI221_X1 port map( B1 => n274, B2 => n2503, C1 => n271, C2 => n3625
                           , A => n1853, ZN => n1858);
   U1512 : OAI22_X1 port map( A1 => n280, A2 => n1855, B1 => n277, B2 => n1854,
                           ZN => n1856);
   U1513 : AOI221_X1 port map( B1 => n286, B2 => n3727, C1 => n283, C2 => n3761
                           , A => n1856, ZN => n1857);
   U1514 : NAND4_X1 port map( A1 => n1860, A2 => n1859, A3 => n1858, A4 => 
                           n1857, ZN => n1861);
   U1515 : OAI21_X1 port map( B1 => n1862, B2 => n1861, A => n289, ZN => n1863)
                           ;
   U1516 : OAI21_X1 port map( B1 => n292, B2 => n1864, A => n1863, ZN => n2581)
                           ;
   U1517 : OAI22_X1 port map( A1 => n196, A2 => n1866, B1 => n193, B2 => n1865,
                           ZN => n1867);
   U1518 : AOI221_X1 port map( B1 => n202, B2 => n3865, C1 => n199, C2 => n3899
                           , A => n1867, ZN => n1880);
   U1519 : OAI22_X1 port map( A1 => n208, A2 => n1869, B1 => n205, B2 => n1868,
                           ZN => n1870);
   U1520 : AOI221_X1 port map( B1 => n214, B2 => n4001, C1 => n211, C2 => n4035
                           , A => n1870, ZN => n1879);
   U1521 : OAI22_X1 port map( A1 => n220, A2 => n1872, B1 => n217, B2 => n1871,
                           ZN => n1873);
   U1522 : AOI221_X1 port map( B1 => n226, B2 => n4141, C1 => n223, C2 => n4176
                           , A => n1873, ZN => n1878);
   U1523 : OAI22_X1 port map( A1 => n232, A2 => n1875, B1 => n229, B2 => n1874,
                           ZN => n1876);
   U1524 : AOI221_X1 port map( B1 => n238, B2 => n4281, C1 => n235, C2 => n4339
                           , A => n1876, ZN => n1877);
   U1525 : NAND4_X1 port map( A1 => n1880, A2 => n1879, A3 => n1878, A4 => 
                           n1877, ZN => n1898);
   U1526 : OAI22_X1 port map( A1 => n244, A2 => n1882, B1 => n241, B2 => n1881,
                           ZN => n1883);
   U1527 : AOI221_X1 port map( B1 => n250, B2 => n2296, C1 => n247, C2 => n2330
                           , A => n1883, ZN => n1896);
   U1528 : OAI22_X1 port map( A1 => n256, A2 => n1885, B1 => n253, B2 => n1884,
                           ZN => n1886);
   U1529 : AOI221_X1 port map( B1 => n262, B2 => n2432, C1 => n259, C2 => n2470
                           , A => n1886, ZN => n1895);
   U1530 : OAI22_X1 port map( A1 => n268, A2 => n1888, B1 => n265, B2 => n1887,
                           ZN => n1889);
   U1531 : AOI221_X1 port map( B1 => n274, B2 => n2504, C1 => n271, C2 => n3626
                           , A => n1889, ZN => n1894);
   U1532 : OAI22_X1 port map( A1 => n280, A2 => n1891, B1 => n277, B2 => n1890,
                           ZN => n1892);
   U1533 : AOI221_X1 port map( B1 => n286, B2 => n3728, C1 => n283, C2 => n3762
                           , A => n1892, ZN => n1893);
   U1534 : NAND4_X1 port map( A1 => n1896, A2 => n1895, A3 => n1894, A4 => 
                           n1893, ZN => n1897);
   U1535 : OAI21_X1 port map( B1 => n1898, B2 => n1897, A => n289, ZN => n1899)
                           ;
   U1536 : OAI21_X1 port map( B1 => n293, B2 => n1900, A => n1899, ZN => n2582)
                           ;
   U1537 : OAI22_X1 port map( A1 => n197, A2 => n1902, B1 => n194, B2 => n1901,
                           ZN => n1903);
   U1538 : AOI221_X1 port map( B1 => n203, B2 => n3866, C1 => n200, C2 => n3900
                           , A => n1903, ZN => n1916);
   U1539 : OAI22_X1 port map( A1 => n209, A2 => n1905, B1 => n206, B2 => n1904,
                           ZN => n1906);
   U1540 : AOI221_X1 port map( B1 => n215, B2 => n4002, C1 => n212, C2 => n4036
                           , A => n1906, ZN => n1915);
   U1541 : OAI22_X1 port map( A1 => n221, A2 => n1908, B1 => n218, B2 => n1907,
                           ZN => n1909);
   U1542 : AOI221_X1 port map( B1 => n227, B2 => n4142, C1 => n224, C2 => n4177
                           , A => n1909, ZN => n1914);
   U1543 : OAI22_X1 port map( A1 => n233, A2 => n1911, B1 => n230, B2 => n1910,
                           ZN => n1912);
   U1544 : AOI221_X1 port map( B1 => n239, B2 => n4282, C1 => n236, C2 => n4341
                           , A => n1912, ZN => n1913);
   U1545 : NAND4_X1 port map( A1 => n1916, A2 => n1915, A3 => n1914, A4 => 
                           n1913, ZN => n1934);
   U1546 : OAI22_X1 port map( A1 => n245, A2 => n1918, B1 => n242, B2 => n1917,
                           ZN => n1919);
   U1547 : AOI221_X1 port map( B1 => n251, B2 => n2297, C1 => n248, C2 => n2331
                           , A => n1919, ZN => n1932);
   U1548 : OAI22_X1 port map( A1 => n257, A2 => n1921, B1 => n254, B2 => n1920,
                           ZN => n1922);
   U1549 : AOI221_X1 port map( B1 => n263, B2 => n2433, C1 => n260, C2 => n2471
                           , A => n1922, ZN => n1931);
   U1550 : OAI22_X1 port map( A1 => n269, A2 => n1924, B1 => n266, B2 => n1923,
                           ZN => n1925);
   U1551 : AOI221_X1 port map( B1 => n275, B2 => n2505, C1 => n272, C2 => n3627
                           , A => n1925, ZN => n1930);
   U1552 : OAI22_X1 port map( A1 => n281, A2 => n1927, B1 => n278, B2 => n1926,
                           ZN => n1928);
   U1553 : AOI221_X1 port map( B1 => n287, B2 => n3729, C1 => n284, C2 => n3763
                           , A => n1928, ZN => n1929);
   U1554 : NAND4_X1 port map( A1 => n1932, A2 => n1931, A3 => n1930, A4 => 
                           n1929, ZN => n1933);
   U1555 : OAI21_X1 port map( B1 => n1934, B2 => n1933, A => n290, ZN => n1935)
                           ;
   U1556 : OAI21_X1 port map( B1 => n293, B2 => n1936, A => n1935, ZN => n2583)
                           ;
   U1557 : OAI22_X1 port map( A1 => n197, A2 => n1938, B1 => n194, B2 => n1937,
                           ZN => n1939);
   U1558 : AOI221_X1 port map( B1 => n203, B2 => n3867, C1 => n200, C2 => n3901
                           , A => n1939, ZN => n1952);
   U1559 : OAI22_X1 port map( A1 => n209, A2 => n1941, B1 => n206, B2 => n1940,
                           ZN => n1942);
   U1560 : AOI221_X1 port map( B1 => n215, B2 => n4003, C1 => n212, C2 => n4037
                           , A => n1942, ZN => n1951);
   U1561 : OAI22_X1 port map( A1 => n221, A2 => n1944, B1 => n218, B2 => n1943,
                           ZN => n1945);
   U1562 : AOI221_X1 port map( B1 => n227, B2 => n4143, C1 => n224, C2 => n4178
                           , A => n1945, ZN => n1950);
   U1563 : OAI22_X1 port map( A1 => n233, A2 => n1947, B1 => n230, B2 => n1946,
                           ZN => n1948);
   U1564 : AOI221_X1 port map( B1 => n239, B2 => n4283, C1 => n236, C2 => n4343
                           , A => n1948, ZN => n1949);
   U1565 : NAND4_X1 port map( A1 => n1952, A2 => n1951, A3 => n1950, A4 => 
                           n1949, ZN => n1970);
   U1566 : OAI22_X1 port map( A1 => n245, A2 => n1954, B1 => n242, B2 => n1953,
                           ZN => n1955);
   U1567 : AOI221_X1 port map( B1 => n251, B2 => n2298, C1 => n248, C2 => n2332
                           , A => n1955, ZN => n1968);
   U1568 : OAI22_X1 port map( A1 => n257, A2 => n1957, B1 => n254, B2 => n1956,
                           ZN => n1958);
   U1569 : AOI221_X1 port map( B1 => n263, B2 => n2434, C1 => n260, C2 => n2472
                           , A => n1958, ZN => n1967);
   U1570 : OAI22_X1 port map( A1 => n269, A2 => n1960, B1 => n266, B2 => n1959,
                           ZN => n1961);
   U1571 : AOI221_X1 port map( B1 => n275, B2 => n2506, C1 => n272, C2 => n3628
                           , A => n1961, ZN => n1966);
   U1572 : OAI22_X1 port map( A1 => n281, A2 => n1963, B1 => n278, B2 => n1962,
                           ZN => n1964);
   U1573 : AOI221_X1 port map( B1 => n287, B2 => n3730, C1 => n284, C2 => n3764
                           , A => n1964, ZN => n1965);
   U1574 : NAND4_X1 port map( A1 => n1968, A2 => n1967, A3 => n1966, A4 => 
                           n1965, ZN => n1969);
   U1575 : OAI21_X1 port map( B1 => n1970, B2 => n1969, A => n290, ZN => n1971)
                           ;
   U1576 : OAI21_X1 port map( B1 => n293, B2 => n6, A => n1971, ZN => n2584);
   U1577 : OAI22_X1 port map( A1 => n197, A2 => n1973, B1 => n194, B2 => n1972,
                           ZN => n1974);
   U1578 : AOI221_X1 port map( B1 => n203, B2 => n3868, C1 => n200, C2 => n3902
                           , A => n1974, ZN => n1987);
   U1579 : OAI22_X1 port map( A1 => n209, A2 => n1976, B1 => n206, B2 => n1975,
                           ZN => n1977);
   U1580 : AOI221_X1 port map( B1 => n215, B2 => n4004, C1 => n212, C2 => n4038
                           , A => n1977, ZN => n1986);
   U1581 : OAI22_X1 port map( A1 => n221, A2 => n1979, B1 => n218, B2 => n1978,
                           ZN => n1980);
   U1582 : AOI221_X1 port map( B1 => n227, B2 => n4144, C1 => n224, C2 => n4179
                           , A => n1980, ZN => n1985);
   U1583 : OAI22_X1 port map( A1 => n233, A2 => n1982, B1 => n230, B2 => n1981,
                           ZN => n1983);
   U1584 : AOI221_X1 port map( B1 => n239, B2 => n4284, C1 => n236, C2 => n4345
                           , A => n1983, ZN => n1984);
   U1585 : NAND4_X1 port map( A1 => n1987, A2 => n1986, A3 => n1985, A4 => 
                           n1984, ZN => n2005);
   U1586 : OAI22_X1 port map( A1 => n245, A2 => n1989, B1 => n242, B2 => n1988,
                           ZN => n1990);
   U1587 : AOI221_X1 port map( B1 => n251, B2 => n2299, C1 => n248, C2 => n2333
                           , A => n1990, ZN => n2003);
   U1588 : OAI22_X1 port map( A1 => n257, A2 => n1992, B1 => n254, B2 => n1991,
                           ZN => n1993);
   U1589 : AOI221_X1 port map( B1 => n263, B2 => n2435, C1 => n260, C2 => n2473
                           , A => n1993, ZN => n2002);
   U1590 : OAI22_X1 port map( A1 => n269, A2 => n1995, B1 => n266, B2 => n1994,
                           ZN => n1996);
   U1591 : AOI221_X1 port map( B1 => n275, B2 => n2507, C1 => n272, C2 => n3629
                           , A => n1996, ZN => n2001);
   U1592 : OAI22_X1 port map( A1 => n281, A2 => n1998, B1 => n278, B2 => n1997,
                           ZN => n1999);
   U1593 : AOI221_X1 port map( B1 => n287, B2 => n3731, C1 => n284, C2 => n3765
                           , A => n1999, ZN => n2000);
   U1594 : NAND4_X1 port map( A1 => n2003, A2 => n2002, A3 => n2001, A4 => 
                           n2000, ZN => n2004);
   U1595 : OAI21_X1 port map( B1 => n2005, B2 => n2004, A => n290, ZN => n2006)
                           ;
   U1596 : OAI21_X1 port map( B1 => n293, B2 => n5, A => n2006, ZN => n2585);
   U1597 : OAI22_X1 port map( A1 => n197, A2 => n2008, B1 => n194, B2 => n2007,
                           ZN => n2009);
   U1598 : AOI221_X1 port map( B1 => n203, B2 => n3869, C1 => n200, C2 => n3903
                           , A => n2009, ZN => n2022);
   U1599 : OAI22_X1 port map( A1 => n209, A2 => n2011, B1 => n206, B2 => n2010,
                           ZN => n2012);
   U1600 : AOI221_X1 port map( B1 => n215, B2 => n4005, C1 => n212, C2 => n4039
                           , A => n2012, ZN => n2021);
   U1601 : OAI22_X1 port map( A1 => n221, A2 => n2014, B1 => n218, B2 => n2013,
                           ZN => n2015);
   U1602 : AOI221_X1 port map( B1 => n227, B2 => n4145, C1 => n224, C2 => n4180
                           , A => n2015, ZN => n2020);
   U1603 : OAI22_X1 port map( A1 => n233, A2 => n2017, B1 => n230, B2 => n2016,
                           ZN => n2018);
   U1604 : AOI221_X1 port map( B1 => n239, B2 => n4285, C1 => n236, C2 => n4347
                           , A => n2018, ZN => n2019);
   U1605 : NAND4_X1 port map( A1 => n2022, A2 => n2021, A3 => n2020, A4 => 
                           n2019, ZN => n2040);
   U1606 : OAI22_X1 port map( A1 => n245, A2 => n2024, B1 => n242, B2 => n2023,
                           ZN => n2025);
   U1607 : AOI221_X1 port map( B1 => n251, B2 => n2300, C1 => n248, C2 => n2334
                           , A => n2025, ZN => n2038);
   U1608 : OAI22_X1 port map( A1 => n257, A2 => n2027, B1 => n254, B2 => n2026,
                           ZN => n2028);
   U1609 : AOI221_X1 port map( B1 => n263, B2 => n2436, C1 => n260, C2 => n2474
                           , A => n2028, ZN => n2037);
   U1610 : OAI22_X1 port map( A1 => n269, A2 => n2030, B1 => n266, B2 => n2029,
                           ZN => n2031);
   U1611 : AOI221_X1 port map( B1 => n275, B2 => n2508, C1 => n272, C2 => n3630
                           , A => n2031, ZN => n2036);
   U1612 : OAI22_X1 port map( A1 => n281, A2 => n2033, B1 => n278, B2 => n2032,
                           ZN => n2034);
   U1613 : AOI221_X1 port map( B1 => n287, B2 => n3732, C1 => n284, C2 => n3766
                           , A => n2034, ZN => n2035);
   U1614 : NAND4_X1 port map( A1 => n2038, A2 => n2037, A3 => n2036, A4 => 
                           n2035, ZN => n2039);
   U1615 : OAI21_X1 port map( B1 => n2040, B2 => n2039, A => n290, ZN => n2041)
                           ;
   U1616 : OAI21_X1 port map( B1 => n293, B2 => n2042, A => n2041, ZN => n2586)
                           ;
   U1617 : OAI22_X1 port map( A1 => n197, A2 => n2044, B1 => n194, B2 => n2043,
                           ZN => n2045);
   U1618 : AOI221_X1 port map( B1 => n203, B2 => n3870, C1 => n200, C2 => n3904
                           , A => n2045, ZN => n2058);
   U1619 : OAI22_X1 port map( A1 => n209, A2 => n2047, B1 => n206, B2 => n2046,
                           ZN => n2048);
   U1620 : AOI221_X1 port map( B1 => n215, B2 => n4006, C1 => n212, C2 => n4040
                           , A => n2048, ZN => n2057);
   U1621 : OAI22_X1 port map( A1 => n221, A2 => n2050, B1 => n218, B2 => n2049,
                           ZN => n2051);
   U1622 : AOI221_X1 port map( B1 => n227, B2 => n4146, C1 => n224, C2 => n4181
                           , A => n2051, ZN => n2056);
   U1623 : OAI22_X1 port map( A1 => n233, A2 => n2053, B1 => n230, B2 => n2052,
                           ZN => n2054);
   U1624 : AOI221_X1 port map( B1 => n239, B2 => n4286, C1 => n236, C2 => n4349
                           , A => n2054, ZN => n2055);
   U1625 : NAND4_X1 port map( A1 => n2058, A2 => n2057, A3 => n2056, A4 => 
                           n2055, ZN => n2076);
   U1626 : OAI22_X1 port map( A1 => n245, A2 => n2060, B1 => n242, B2 => n2059,
                           ZN => n2061);
   U1627 : AOI221_X1 port map( B1 => n251, B2 => n2301, C1 => n248, C2 => n2335
                           , A => n2061, ZN => n2074);
   U1628 : OAI22_X1 port map( A1 => n257, A2 => n2063, B1 => n254, B2 => n2062,
                           ZN => n2064);
   U1629 : AOI221_X1 port map( B1 => n263, B2 => n2437, C1 => n260, C2 => n2475
                           , A => n2064, ZN => n2073);
   U1630 : OAI22_X1 port map( A1 => n269, A2 => n2066, B1 => n266, B2 => n2065,
                           ZN => n2067);
   U1631 : AOI221_X1 port map( B1 => n275, B2 => n2509, C1 => n272, C2 => n3631
                           , A => n2067, ZN => n2072);
   U1632 : OAI22_X1 port map( A1 => n281, A2 => n2069, B1 => n278, B2 => n2068,
                           ZN => n2070);
   U1633 : AOI221_X1 port map( B1 => n287, B2 => n3733, C1 => n284, C2 => n3767
                           , A => n2070, ZN => n2071);
   U1634 : NAND4_X1 port map( A1 => n2074, A2 => n2073, A3 => n2072, A4 => 
                           n2071, ZN => n2075);
   U1635 : OAI21_X1 port map( B1 => n2076, B2 => n2075, A => n290, ZN => n2077)
                           ;
   U1636 : OAI21_X1 port map( B1 => n293, B2 => n2078, A => n2077, ZN => n2587)
                           ;
   U1637 : OAI22_X1 port map( A1 => n197, A2 => n2080, B1 => n194, B2 => n2079,
                           ZN => n2081);
   U1638 : AOI221_X1 port map( B1 => n203, B2 => n3871, C1 => n200, C2 => n3905
                           , A => n2081, ZN => n2094);
   U1639 : OAI22_X1 port map( A1 => n209, A2 => n2083, B1 => n206, B2 => n2082,
                           ZN => n2084);
   U1640 : AOI221_X1 port map( B1 => n215, B2 => n4007, C1 => n212, C2 => n4041
                           , A => n2084, ZN => n2093);
   U1641 : OAI22_X1 port map( A1 => n221, A2 => n2086, B1 => n218, B2 => n2085,
                           ZN => n2087);
   U1642 : AOI221_X1 port map( B1 => n227, B2 => n4147, C1 => n224, C2 => n4182
                           , A => n2087, ZN => n2092);
   U1643 : OAI22_X1 port map( A1 => n233, A2 => n2089, B1 => n230, B2 => n2088,
                           ZN => n2090);
   U1644 : AOI221_X1 port map( B1 => n239, B2 => n4287, C1 => n236, C2 => n4351
                           , A => n2090, ZN => n2091);
   U1645 : NAND4_X1 port map( A1 => n2094, A2 => n2093, A3 => n2092, A4 => 
                           n2091, ZN => n2112);
   U1646 : OAI22_X1 port map( A1 => n245, A2 => n2096, B1 => n242, B2 => n2095,
                           ZN => n2097);
   U1647 : AOI221_X1 port map( B1 => n251, B2 => n2302, C1 => n248, C2 => n2336
                           , A => n2097, ZN => n2110);
   U1648 : OAI22_X1 port map( A1 => n257, A2 => n2099, B1 => n254, B2 => n2098,
                           ZN => n2100);
   U1649 : AOI221_X1 port map( B1 => n263, B2 => n2438, C1 => n260, C2 => n2476
                           , A => n2100, ZN => n2109);
   U1650 : OAI22_X1 port map( A1 => n269, A2 => n2102, B1 => n266, B2 => n2101,
                           ZN => n2103);
   U1651 : AOI221_X1 port map( B1 => n275, B2 => n2510, C1 => n272, C2 => n3632
                           , A => n2103, ZN => n2108);
   U1652 : OAI22_X1 port map( A1 => n281, A2 => n2105, B1 => n278, B2 => n2104,
                           ZN => n2106);
   U1653 : AOI221_X1 port map( B1 => n287, B2 => n3734, C1 => n284, C2 => n3768
                           , A => n2106, ZN => n2107);
   U1654 : NAND4_X1 port map( A1 => n2110, A2 => n2109, A3 => n2108, A4 => 
                           n2107, ZN => n2111);
   U1655 : OAI21_X1 port map( B1 => n2112, B2 => n2111, A => n290, ZN => n2113)
                           ;
   U1656 : OAI21_X1 port map( B1 => n293, B2 => n2114, A => n2113, ZN => n2588)
                           ;
   U1657 : OAI22_X1 port map( A1 => n197, A2 => n2116, B1 => n194, B2 => n2115,
                           ZN => n2117);
   U1658 : AOI221_X1 port map( B1 => n203, B2 => n3872, C1 => n200, C2 => n3906
                           , A => n2117, ZN => n2130);
   U1659 : OAI22_X1 port map( A1 => n209, A2 => n2119, B1 => n206, B2 => n2118,
                           ZN => n2120);
   U1660 : AOI221_X1 port map( B1 => n215, B2 => n4008, C1 => n212, C2 => n4042
                           , A => n2120, ZN => n2129);
   U1661 : OAI22_X1 port map( A1 => n221, A2 => n2122, B1 => n218, B2 => n2121,
                           ZN => n2123);
   U1662 : AOI221_X1 port map( B1 => n227, B2 => n4148, C1 => n224, C2 => n4183
                           , A => n2123, ZN => n2128);
   U1663 : OAI22_X1 port map( A1 => n233, A2 => n2125, B1 => n230, B2 => n2124,
                           ZN => n2126);
   U1664 : AOI221_X1 port map( B1 => n239, B2 => n4288, C1 => n236, C2 => n4353
                           , A => n2126, ZN => n2127);
   U1665 : NAND4_X1 port map( A1 => n2130, A2 => n2129, A3 => n2128, A4 => 
                           n2127, ZN => n2148);
   U1666 : OAI22_X1 port map( A1 => n245, A2 => n2132, B1 => n242, B2 => n2131,
                           ZN => n2133);
   U1667 : AOI221_X1 port map( B1 => n251, B2 => n2303, C1 => n248, C2 => n2337
                           , A => n2133, ZN => n2146);
   U1668 : OAI22_X1 port map( A1 => n257, A2 => n2135, B1 => n254, B2 => n2134,
                           ZN => n2136);
   U1669 : AOI221_X1 port map( B1 => n263, B2 => n2439, C1 => n260, C2 => n2477
                           , A => n2136, ZN => n2145);
   U1670 : OAI22_X1 port map( A1 => n269, A2 => n2138, B1 => n266, B2 => n2137,
                           ZN => n2139);
   U1671 : AOI221_X1 port map( B1 => n275, B2 => n2511, C1 => n272, C2 => n3633
                           , A => n2139, ZN => n2144);
   U1672 : OAI22_X1 port map( A1 => n281, A2 => n2141, B1 => n278, B2 => n2140,
                           ZN => n2142);
   U1673 : AOI221_X1 port map( B1 => n287, B2 => n3735, C1 => n284, C2 => n3769
                           , A => n2142, ZN => n2143);
   U1674 : NAND4_X1 port map( A1 => n2146, A2 => n2145, A3 => n2144, A4 => 
                           n2143, ZN => n2147);
   U1675 : OAI21_X1 port map( B1 => n2148, B2 => n2147, A => n290, ZN => n2149)
                           ;
   U1676 : OAI21_X1 port map( B1 => n293, B2 => n2150, A => n2149, ZN => n2589)
                           ;
   U1677 : OAI22_X1 port map( A1 => n197, A2 => n2153, B1 => n194, B2 => n2151,
                           ZN => n2155);
   U1678 : AOI221_X1 port map( B1 => n203, B2 => n3874, C1 => n200, C2 => n3908
                           , A => n2155, ZN => n2174);
   U1679 : OAI22_X1 port map( A1 => n209, A2 => n2158, B1 => n206, B2 => n2156,
                           ZN => n2160);
   U1680 : AOI221_X1 port map( B1 => n215, B2 => n4010, C1 => n212, C2 => n4044
                           , A => n2160, ZN => n2173);
   U1681 : OAI22_X1 port map( A1 => n221, A2 => n2163, B1 => n218, B2 => n2161,
                           ZN => n2165);
   U1682 : AOI221_X1 port map( B1 => n227, B2 => n4150, C1 => n224, C2 => n4185
                           , A => n2165, ZN => n2172);
   U1683 : OAI22_X1 port map( A1 => n233, A2 => n2168, B1 => n230, B2 => n2166,
                           ZN => n2170);
   U1684 : AOI221_X1 port map( B1 => n239, B2 => n4290, C1 => n236, C2 => n4356
                           , A => n2170, ZN => n2171);
   U1685 : NAND4_X1 port map( A1 => n2174, A2 => n2173, A3 => n2172, A4 => 
                           n2171, ZN => n2200);
   U1686 : OAI22_X1 port map( A1 => n245, A2 => n2177, B1 => n242, B2 => n2175,
                           ZN => n2179);
   U1687 : AOI221_X1 port map( B1 => n251, B2 => n2305, C1 => n248, C2 => n2339
                           , A => n2179, ZN => n2198);
   U1688 : OAI22_X1 port map( A1 => n257, A2 => n2182, B1 => n254, B2 => n2180,
                           ZN => n2184);
   U1689 : AOI221_X1 port map( B1 => n263, B2 => n2441, C1 => n260, C2 => n2479
                           , A => n2184, ZN => n2197);
   U1690 : OAI22_X1 port map( A1 => n269, A2 => n2187, B1 => n266, B2 => n2185,
                           ZN => n2189);
   U1691 : AOI221_X1 port map( B1 => n275, B2 => n2513, C1 => n272, C2 => n3635
                           , A => n2189, ZN => n2196);
   U1692 : OAI22_X1 port map( A1 => n281, A2 => n2192, B1 => n278, B2 => n2190,
                           ZN => n2194);
   U1693 : AOI221_X1 port map( B1 => n287, B2 => n3737, C1 => n284, C2 => n3771
                           , A => n2194, ZN => n2195);
   U1694 : NAND4_X1 port map( A1 => n2198, A2 => n2197, A3 => n2196, A4 => 
                           n2195, ZN => n2199);
   U1695 : OAI21_X1 port map( B1 => n2200, B2 => n2199, A => n290, ZN => n2201)
                           ;
   U1696 : OAI21_X1 port map( B1 => n293, B2 => n2202, A => n2201, ZN => n2590)
                           ;
   U1697 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n85, ZN => n4396);
   U1698 : NAND2_X1 port map( A1 => n15, A2 => ADD_WR(0), ZN => n4116);
   U1699 : NAND2_X1 port map( A1 => n16, A2 => ADD_WR(3), ZN => n2445);
   U1700 : OAI21_X1 port map( B1 => n4116, B2 => n2445, A => n83, ZN => n2204);
   U1701 : INV_X1 port map( A => n2204, ZN => n2236);
   U1702 : MUX2_X1 port map( A => n4396, B => n1060, S => n294, Z => n2205);
   U1703 : INV_X1 port map( A => n2205, ZN => n2591);
   U1704 : MUX2_X1 port map( A => n4398, B => n1098, S => n294, Z => n2206);
   U1705 : INV_X1 port map( A => n2206, ZN => n2592);
   U1706 : MUX2_X1 port map( A => n4400, B => n1134, S => n294, Z => n2207);
   U1707 : INV_X1 port map( A => n2207, ZN => n2593);
   U1708 : MUX2_X1 port map( A => n4402, B => n1170, S => n294, Z => n2208);
   U1709 : INV_X1 port map( A => n2208, ZN => n2594);
   U1710 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n85, ZN => n4404);
   U1711 : MUX2_X1 port map( A => n4404, B => n1206, S => n294, Z => n2209);
   U1712 : INV_X1 port map( A => n2209, ZN => n2595);
   U1713 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n83, ZN => n4406);
   U1714 : MUX2_X1 port map( A => n4406, B => n1242, S => n294, Z => n2210);
   U1715 : INV_X1 port map( A => n2210, ZN => n2596);
   U1716 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n85, ZN => n4408);
   U1717 : MUX2_X1 port map( A => n4408, B => n1278, S => n294, Z => n2211);
   U1718 : INV_X1 port map( A => n2211, ZN => n2597);
   U1719 : NAND2_X1 port map( A1 => DATAIN(7), A2 => RST, ZN => n4410);
   U1720 : MUX2_X1 port map( A => n4410, B => n1314, S => n294, Z => n2212);
   U1721 : INV_X1 port map( A => n2212, ZN => n2598);
   U1722 : NAND2_X1 port map( A1 => DATAIN(8), A2 => RST, ZN => n4412);
   U1723 : MUX2_X1 port map( A => n4412, B => n1350, S => n294, Z => n2213);
   U1724 : INV_X1 port map( A => n2213, ZN => n2599);
   U1725 : NAND2_X1 port map( A1 => DATAIN(9), A2 => RST, ZN => n4414);
   U1726 : MUX2_X1 port map( A => n4414, B => n1385, S => n294, Z => n2214);
   U1727 : INV_X1 port map( A => n2214, ZN => n2600);
   U1728 : NAND2_X1 port map( A1 => DATAIN(10), A2 => RST, ZN => n4416);
   U1729 : MUX2_X1 port map( A => n4416, B => n1420, S => n294, Z => n2215);
   U1730 : INV_X1 port map( A => n2215, ZN => n2601);
   U1731 : NAND2_X1 port map( A1 => DATAIN(11), A2 => RST, ZN => n4418);
   U1732 : MUX2_X1 port map( A => n4418, B => n1455, S => n294, Z => n2216);
   U1733 : INV_X1 port map( A => n2216, ZN => n2602);
   U1734 : NAND2_X1 port map( A1 => DATAIN(12), A2 => RST, ZN => n4420);
   U1735 : MUX2_X1 port map( A => n4420, B => n1490, S => n295, Z => n2217);
   U1736 : INV_X1 port map( A => n2217, ZN => n2603);
   U1737 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n85, ZN => n4422);
   U1738 : MUX2_X1 port map( A => n4422, B => n1525, S => n295, Z => n2218);
   U1739 : INV_X1 port map( A => n2218, ZN => n2604);
   U1740 : NAND2_X1 port map( A1 => DATAIN(14), A2 => RST, ZN => n4424);
   U1741 : MUX2_X1 port map( A => n4424, B => n1561, S => n295, Z => n2219);
   U1742 : INV_X1 port map( A => n2219, ZN => n2605);
   U1743 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n84, ZN => n4426);
   U1744 : MUX2_X1 port map( A => n4426, B => n1596, S => n295, Z => n2220);
   U1745 : INV_X1 port map( A => n2220, ZN => n2606);
   U1746 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n84, ZN => n4428);
   U1747 : MUX2_X1 port map( A => n4428, B => n1631, S => n295, Z => n2221);
   U1748 : INV_X1 port map( A => n2221, ZN => n2607);
   U1749 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n85, ZN => n4430);
   U1750 : MUX2_X1 port map( A => n4430, B => n1667, S => n295, Z => n2222);
   U1751 : INV_X1 port map( A => n2222, ZN => n2608);
   U1752 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n85, ZN => n4432);
   U1753 : MUX2_X1 port map( A => n4432, B => n1703, S => n295, Z => n2223);
   U1754 : INV_X1 port map( A => n2223, ZN => n2609);
   U1755 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n85, ZN => n4434);
   U1756 : MUX2_X1 port map( A => n4434, B => n1738, S => n295, Z => n2224);
   U1757 : INV_X1 port map( A => n2224, ZN => n2610);
   U1758 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n85, ZN => n4436);
   U1759 : MUX2_X1 port map( A => n4436, B => n1774, S => n295, Z => n2225);
   U1760 : INV_X1 port map( A => n2225, ZN => n2611);
   U1761 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n85, ZN => n4438);
   U1762 : MUX2_X1 port map( A => n4438, B => n1810, S => n295, Z => n2226);
   U1763 : INV_X1 port map( A => n2226, ZN => n2612);
   U1764 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n85, ZN => n4440);
   U1765 : MUX2_X1 port map( A => n4440, B => n1846, S => n295, Z => n2227);
   U1766 : INV_X1 port map( A => n2227, ZN => n2613);
   U1767 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n85, ZN => n4442);
   U1768 : MUX2_X1 port map( A => n4442, B => n1882, S => n295, Z => n2228);
   U1769 : INV_X1 port map( A => n2228, ZN => n2614);
   U1770 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n85, ZN => n4444);
   U1771 : MUX2_X1 port map( A => n4444, B => n1918, S => n296, Z => n2229);
   U1772 : INV_X1 port map( A => n2229, ZN => n2615);
   U1773 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n85, ZN => n4446);
   U1774 : MUX2_X1 port map( A => n4446, B => n1954, S => n296, Z => n2230);
   U1775 : INV_X1 port map( A => n2230, ZN => n2616);
   U1776 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n85, ZN => n4448);
   U1777 : MUX2_X1 port map( A => n4448, B => n1989, S => n296, Z => n2231);
   U1778 : INV_X1 port map( A => n2231, ZN => n2617);
   U1779 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n85, ZN => n4450);
   U1780 : MUX2_X1 port map( A => n4450, B => n2024, S => n296, Z => n2232);
   U1781 : INV_X1 port map( A => n2232, ZN => n2618);
   U1782 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n85, ZN => n4452);
   U1783 : MUX2_X1 port map( A => n4452, B => n2060, S => n296, Z => n2233);
   U1784 : INV_X1 port map( A => n2233, ZN => n2619);
   U1785 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n84, ZN => n4454);
   U1786 : MUX2_X1 port map( A => n4454, B => n2096, S => n296, Z => n2234);
   U1787 : INV_X1 port map( A => n2234, ZN => n2620);
   U1788 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n85, ZN => n4456);
   U1789 : MUX2_X1 port map( A => n4456, B => n2132, S => n296, Z => n2235);
   U1790 : INV_X1 port map( A => n2235, ZN => n2621);
   U1791 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n85, ZN => n4459);
   U1792 : MUX2_X1 port map( A => n4459, B => n2177, S => n296, Z => n2237);
   U1793 : INV_X1 port map( A => n2237, ZN => n2622);
   U1794 : INV_X1 port map( A => ADD_WR(0), ZN => n2442);
   U1795 : NAND2_X1 port map( A1 => n15, A2 => n2442, ZN => n4151);
   U1796 : OAI21_X1 port map( B1 => n4151, B2 => n2445, A => n84, ZN => n2238);
   U1797 : INV_X1 port map( A => n2238, ZN => n2270);
   U1798 : MUX2_X1 port map( A => n4396, B => n1059, S => n297, Z => n2239);
   U1799 : INV_X1 port map( A => n2239, ZN => n2623);
   U1800 : MUX2_X1 port map( A => n4398, B => n1097, S => n297, Z => n2240);
   U1801 : INV_X1 port map( A => n2240, ZN => n2624);
   U1802 : MUX2_X1 port map( A => n4400, B => n1133, S => n297, Z => n2241);
   U1803 : INV_X1 port map( A => n2241, ZN => n2625);
   U1804 : MUX2_X1 port map( A => n4402, B => n1169, S => n297, Z => n2242);
   U1805 : INV_X1 port map( A => n2242, ZN => n2626);
   U1806 : MUX2_X1 port map( A => n4404, B => n1205, S => n297, Z => n2243);
   U1807 : INV_X1 port map( A => n2243, ZN => n2627);
   U1808 : MUX2_X1 port map( A => n4406, B => n1241, S => n297, Z => n2244);
   U1809 : INV_X1 port map( A => n2244, ZN => n2628);
   U1810 : MUX2_X1 port map( A => n4408, B => n1277, S => n297, Z => n2245);
   U1811 : INV_X1 port map( A => n2245, ZN => n2629);
   U1812 : MUX2_X1 port map( A => n4410, B => n1313, S => n297, Z => n2246);
   U1813 : INV_X1 port map( A => n2246, ZN => n2630);
   U1814 : MUX2_X1 port map( A => n4412, B => n1349, S => n297, Z => n2247);
   U1815 : INV_X1 port map( A => n2247, ZN => n2631);
   U1816 : MUX2_X1 port map( A => n4414, B => n1384, S => n297, Z => n2248);
   U1817 : INV_X1 port map( A => n2248, ZN => n2632);
   U1818 : MUX2_X1 port map( A => n4416, B => n1419, S => n297, Z => n2249);
   U1819 : INV_X1 port map( A => n2249, ZN => n2633);
   U1820 : MUX2_X1 port map( A => n4418, B => n1454, S => n297, Z => n2250);
   U1821 : INV_X1 port map( A => n2250, ZN => n2634);
   U1822 : MUX2_X1 port map( A => n4420, B => n1489, S => n298, Z => n2251);
   U1823 : INV_X1 port map( A => n2251, ZN => n2635);
   U1824 : MUX2_X1 port map( A => n4422, B => n1524, S => n298, Z => n2252);
   U1825 : INV_X1 port map( A => n2252, ZN => n2636);
   U1826 : MUX2_X1 port map( A => n4424, B => n1560, S => n298, Z => n2253);
   U1827 : INV_X1 port map( A => n2253, ZN => n2637);
   U1828 : MUX2_X1 port map( A => n4426, B => n1595, S => n298, Z => n2254);
   U1829 : INV_X1 port map( A => n2254, ZN => n2638);
   U1830 : MUX2_X1 port map( A => n4428, B => n1630, S => n298, Z => n2255);
   U1831 : INV_X1 port map( A => n2255, ZN => n2639);
   U1832 : MUX2_X1 port map( A => n4430, B => n1666, S => n298, Z => n2256);
   U1833 : INV_X1 port map( A => n2256, ZN => n2640);
   U1834 : MUX2_X1 port map( A => n4432, B => n1702, S => n298, Z => n2257);
   U1835 : INV_X1 port map( A => n2257, ZN => n2641);
   U1836 : MUX2_X1 port map( A => n4434, B => n1737, S => n298, Z => n2258);
   U1837 : INV_X1 port map( A => n2258, ZN => n2642);
   U1838 : MUX2_X1 port map( A => n4436, B => n1773, S => n298, Z => n2259);
   U1839 : INV_X1 port map( A => n2259, ZN => n2643);
   U1840 : MUX2_X1 port map( A => n4438, B => n1809, S => n298, Z => n2260);
   U1841 : INV_X1 port map( A => n2260, ZN => n2644);
   U1842 : MUX2_X1 port map( A => n4440, B => n1845, S => n298, Z => n2261);
   U1843 : INV_X1 port map( A => n2261, ZN => n2645);
   U1844 : MUX2_X1 port map( A => n4442, B => n1881, S => n298, Z => n2262);
   U1845 : INV_X1 port map( A => n2262, ZN => n2646);
   U1846 : MUX2_X1 port map( A => n4444, B => n1917, S => n299, Z => n2263);
   U1847 : INV_X1 port map( A => n2263, ZN => n2647);
   U1848 : MUX2_X1 port map( A => n4446, B => n1953, S => n299, Z => n2264);
   U1849 : INV_X1 port map( A => n2264, ZN => n2648);
   U1850 : MUX2_X1 port map( A => n4448, B => n1988, S => n299, Z => n2265);
   U1851 : INV_X1 port map( A => n2265, ZN => n2649);
   U1852 : MUX2_X1 port map( A => n4450, B => n2023, S => n299, Z => n2266);
   U1853 : INV_X1 port map( A => n2266, ZN => n2650);
   U1854 : MUX2_X1 port map( A => n4452, B => n2059, S => n299, Z => n2267);
   U1855 : INV_X1 port map( A => n2267, ZN => n2651);
   U1856 : MUX2_X1 port map( A => n4454, B => n2095, S => n299, Z => n2268);
   U1857 : INV_X1 port map( A => n2268, ZN => n2652);
   U1858 : MUX2_X1 port map( A => n4456, B => n2131, S => n299, Z => n2269);
   U1859 : INV_X1 port map( A => n2269, ZN => n2653);
   U1860 : MUX2_X1 port map( A => n4459, B => n2175, S => n299, Z => n2271);
   U1861 : INV_X1 port map( A => n2271, ZN => n2654);
   U1862 : INV_X1 port map( A => n4396, ZN => n4294);
   U1863 : INV_X1 port map( A => ADD_WR(1), ZN => n2443);
   U1864 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => n2443, ZN
                           => n4186);
   U1865 : OAI21_X1 port map( B1 => n4186, B2 => n2445, A => n84, ZN => n2272);
   U1866 : INV_X1 port map( A => n2272, ZN => n2304);
   U1867 : MUX2_X1 port map( A => n4294, B => n2273, S => n300, Z => n2655);
   U1868 : INV_X1 port map( A => n4398, ZN => n4296);
   U1869 : MUX2_X1 port map( A => n4296, B => n2274, S => n300, Z => n2656);
   U1870 : INV_X1 port map( A => n4400, ZN => n4298);
   U1871 : MUX2_X1 port map( A => n4298, B => n2275, S => n300, Z => n2657);
   U1872 : INV_X1 port map( A => n4402, ZN => n4300);
   U1873 : MUX2_X1 port map( A => n4300, B => n2276, S => n300, Z => n2658);
   U1874 : INV_X1 port map( A => n4404, ZN => n4302);
   U1875 : MUX2_X1 port map( A => n4302, B => n2277, S => n300, Z => n2659);
   U1876 : INV_X1 port map( A => n4406, ZN => n4304);
   U1877 : MUX2_X1 port map( A => n4304, B => n2278, S => n300, Z => n2660);
   U1878 : INV_X1 port map( A => n4408, ZN => n4306);
   U1879 : MUX2_X1 port map( A => n4306, B => n2279, S => n300, Z => n2661);
   U1880 : INV_X1 port map( A => n4410, ZN => n4308);
   U1881 : MUX2_X1 port map( A => n4308, B => n2280, S => n300, Z => n2662);
   U1882 : INV_X1 port map( A => n4412, ZN => n4310);
   U1883 : MUX2_X1 port map( A => n4310, B => n2281, S => n300, Z => n2663);
   U1884 : INV_X1 port map( A => n4414, ZN => n4312);
   U1885 : MUX2_X1 port map( A => n4312, B => n2282, S => n300, Z => n2664);
   U1886 : INV_X1 port map( A => n4416, ZN => n4314);
   U1887 : MUX2_X1 port map( A => n4314, B => n2283, S => n300, Z => n2665);
   U1888 : INV_X1 port map( A => n4418, ZN => n4316);
   U1889 : MUX2_X1 port map( A => n4316, B => n2284, S => n300, Z => n2666);
   U1890 : INV_X1 port map( A => n4420, ZN => n4318);
   U1891 : MUX2_X1 port map( A => n4318, B => n2285, S => n301, Z => n2667);
   U1892 : INV_X1 port map( A => n4422, ZN => n4320);
   U1893 : MUX2_X1 port map( A => n4320, B => n2286, S => n301, Z => n2668);
   U1894 : INV_X1 port map( A => n4424, ZN => n4322);
   U1895 : MUX2_X1 port map( A => n4322, B => n2287, S => n301, Z => n2669);
   U1896 : INV_X1 port map( A => n4426, ZN => n4324);
   U1897 : MUX2_X1 port map( A => n4324, B => n2288, S => n301, Z => n2670);
   U1898 : INV_X1 port map( A => n4428, ZN => n4326);
   U1899 : MUX2_X1 port map( A => n4326, B => n2289, S => n301, Z => n2671);
   U1900 : INV_X1 port map( A => n4430, ZN => n4328);
   U1901 : MUX2_X1 port map( A => n4328, B => n2290, S => n301, Z => n2672);
   U1902 : INV_X1 port map( A => n4432, ZN => n4330);
   U1903 : MUX2_X1 port map( A => n4330, B => n2291, S => n301, Z => n2673);
   U1904 : INV_X1 port map( A => n4434, ZN => n4332);
   U1905 : MUX2_X1 port map( A => n4332, B => n2292, S => n301, Z => n2674);
   U1906 : INV_X1 port map( A => n4436, ZN => n4334);
   U1907 : MUX2_X1 port map( A => n4334, B => n2293, S => n301, Z => n2675);
   U1908 : INV_X1 port map( A => n4438, ZN => n4336);
   U1909 : MUX2_X1 port map( A => n4336, B => n2294, S => n301, Z => n2676);
   U1910 : INV_X1 port map( A => n4440, ZN => n4338);
   U1911 : MUX2_X1 port map( A => n4338, B => n2295, S => n301, Z => n2677);
   U1912 : INV_X1 port map( A => n4442, ZN => n4340);
   U1913 : MUX2_X1 port map( A => n4340, B => n2296, S => n301, Z => n2678);
   U1914 : INV_X1 port map( A => n4444, ZN => n4342);
   U1915 : MUX2_X1 port map( A => n4342, B => n2297, S => n302, Z => n2679);
   U1916 : INV_X1 port map( A => n4446, ZN => n4344);
   U1917 : MUX2_X1 port map( A => n4344, B => n2298, S => n302, Z => n2680);
   U1918 : INV_X1 port map( A => n4448, ZN => n4346);
   U1919 : MUX2_X1 port map( A => n4346, B => n2299, S => n302, Z => n2681);
   U1920 : INV_X1 port map( A => n4450, ZN => n4348);
   U1921 : MUX2_X1 port map( A => n4348, B => n2300, S => n302, Z => n2682);
   U1922 : INV_X1 port map( A => n4452, ZN => n4350);
   U1923 : MUX2_X1 port map( A => n4350, B => n2301, S => n302, Z => n2683);
   U1924 : INV_X1 port map( A => n4454, ZN => n4352);
   U1925 : MUX2_X1 port map( A => n4352, B => n2302, S => n302, Z => n2684);
   U1926 : INV_X1 port map( A => n4456, ZN => n4354);
   U1927 : MUX2_X1 port map( A => n4354, B => n2303, S => n302, Z => n2685);
   U1928 : INV_X1 port map( A => n4459, ZN => n4357);
   U1929 : MUX2_X1 port map( A => n4357, B => n2305, S => n302, Z => n2686);
   U1930 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n2443, A3 => n2442, ZN => 
                           n4221);
   U1931 : OAI21_X1 port map( B1 => n4221, B2 => n2445, A => n84, ZN => n2306);
   U1932 : INV_X1 port map( A => n2306, ZN => n2338);
   U1933 : MUX2_X1 port map( A => n4294, B => n2307, S => n303, Z => n2687);
   U1934 : MUX2_X1 port map( A => n4296, B => n2308, S => n303, Z => n2688);
   U1935 : MUX2_X1 port map( A => n4298, B => n2309, S => n303, Z => n2689);
   U1936 : MUX2_X1 port map( A => n4300, B => n2310, S => n303, Z => n2690);
   U1937 : MUX2_X1 port map( A => n4302, B => n2311, S => n303, Z => n2691);
   U1938 : MUX2_X1 port map( A => n4304, B => n2312, S => n303, Z => n2692);
   U1939 : MUX2_X1 port map( A => n4306, B => n2313, S => n303, Z => n2693);
   U1940 : MUX2_X1 port map( A => n4308, B => n2314, S => n303, Z => n2694);
   U1941 : MUX2_X1 port map( A => n4310, B => n2315, S => n303, Z => n2695);
   U1942 : MUX2_X1 port map( A => n4312, B => n2316, S => n303, Z => n2696);
   U1943 : MUX2_X1 port map( A => n4314, B => n2317, S => n303, Z => n2697);
   U1944 : MUX2_X1 port map( A => n4316, B => n2318, S => n303, Z => n2698);
   U1945 : MUX2_X1 port map( A => n4318, B => n2319, S => n304, Z => n2699);
   U1946 : MUX2_X1 port map( A => n4320, B => n2320, S => n304, Z => n2700);
   U1947 : MUX2_X1 port map( A => n4322, B => n2321, S => n304, Z => n2701);
   U1948 : MUX2_X1 port map( A => n4324, B => n2322, S => n304, Z => n2702);
   U1949 : MUX2_X1 port map( A => n4326, B => n2323, S => n304, Z => n2703);
   U1950 : MUX2_X1 port map( A => n4328, B => n2324, S => n304, Z => n2704);
   U1951 : MUX2_X1 port map( A => n4330, B => n2325, S => n304, Z => n2705);
   U1952 : MUX2_X1 port map( A => n4332, B => n2326, S => n304, Z => n2706);
   U1953 : MUX2_X1 port map( A => n4334, B => n2327, S => n304, Z => n2707);
   U1954 : MUX2_X1 port map( A => n4336, B => n2328, S => n304, Z => n2708);
   U1955 : MUX2_X1 port map( A => n4338, B => n2329, S => n304, Z => n2709);
   U1956 : MUX2_X1 port map( A => n4340, B => n2330, S => n304, Z => n2710);
   U1957 : MUX2_X1 port map( A => n4342, B => n2331, S => n305, Z => n2711);
   U1958 : MUX2_X1 port map( A => n4344, B => n2332, S => n305, Z => n2712);
   U1959 : MUX2_X1 port map( A => n4346, B => n2333, S => n305, Z => n2713);
   U1960 : MUX2_X1 port map( A => n4348, B => n2334, S => n305, Z => n2714);
   U1961 : MUX2_X1 port map( A => n4350, B => n2335, S => n305, Z => n2715);
   U1962 : MUX2_X1 port map( A => n4352, B => n2336, S => n305, Z => n2716);
   U1963 : MUX2_X1 port map( A => n4354, B => n2337, S => n305, Z => n2717);
   U1964 : MUX2_X1 port map( A => n4357, B => n2339, S => n305, Z => n2718);
   U1965 : INV_X1 port map( A => ADD_WR(2), ZN => n2444);
   U1966 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => n2444, ZN
                           => n4256);
   U1967 : OAI21_X1 port map( B1 => n4256, B2 => n2445, A => n84, ZN => n2340);
   U1968 : INV_X1 port map( A => n2340, ZN => n2372);
   U1969 : MUX2_X1 port map( A => n4396, B => n1063, S => n306, Z => n2341);
   U1970 : INV_X1 port map( A => n2341, ZN => n2719);
   U1971 : MUX2_X1 port map( A => n4398, B => n1101, S => n306, Z => n2342);
   U1972 : INV_X1 port map( A => n2342, ZN => n2720);
   U1973 : MUX2_X1 port map( A => n4400, B => n1137, S => n306, Z => n2343);
   U1974 : INV_X1 port map( A => n2343, ZN => n2721);
   U1975 : MUX2_X1 port map( A => n4402, B => n1173, S => n306, Z => n2344);
   U1976 : INV_X1 port map( A => n2344, ZN => n2722);
   U1977 : MUX2_X1 port map( A => n4404, B => n1209, S => n306, Z => n2345);
   U1978 : INV_X1 port map( A => n2345, ZN => n2723);
   U1979 : MUX2_X1 port map( A => n4406, B => n1245, S => n306, Z => n2346);
   U1980 : INV_X1 port map( A => n2346, ZN => n2724);
   U1981 : MUX2_X1 port map( A => n4408, B => n1281, S => n306, Z => n2347);
   U1982 : INV_X1 port map( A => n2347, ZN => n2725);
   U1983 : MUX2_X1 port map( A => n4410, B => n1317, S => n306, Z => n2348);
   U1984 : INV_X1 port map( A => n2348, ZN => n2726);
   U1985 : MUX2_X1 port map( A => n4412, B => n1353, S => n306, Z => n2349);
   U1986 : INV_X1 port map( A => n2349, ZN => n2727);
   U1987 : MUX2_X1 port map( A => n4414, B => n1388, S => n306, Z => n2350);
   U1988 : INV_X1 port map( A => n2350, ZN => n2728);
   U1989 : MUX2_X1 port map( A => n4416, B => n1423, S => n306, Z => n2351);
   U1990 : INV_X1 port map( A => n2351, ZN => n2729);
   U1991 : MUX2_X1 port map( A => n4418, B => n1458, S => n306, Z => n2352);
   U1992 : INV_X1 port map( A => n2352, ZN => n2730);
   U1993 : MUX2_X1 port map( A => n4420, B => n1493, S => n307, Z => n2353);
   U1994 : INV_X1 port map( A => n2353, ZN => n2731);
   U1995 : MUX2_X1 port map( A => n4422, B => n1528, S => n307, Z => n2354);
   U1996 : INV_X1 port map( A => n2354, ZN => n2732);
   U1997 : MUX2_X1 port map( A => n4424, B => n1564, S => n307, Z => n2355);
   U1998 : INV_X1 port map( A => n2355, ZN => n2733);
   U1999 : MUX2_X1 port map( A => n4426, B => n1599, S => n307, Z => n2356);
   U2000 : INV_X1 port map( A => n2356, ZN => n2734);
   U2001 : MUX2_X1 port map( A => n4428, B => n1634, S => n307, Z => n2357);
   U2002 : INV_X1 port map( A => n2357, ZN => n2735);
   U2003 : MUX2_X1 port map( A => n4430, B => n1670, S => n307, Z => n2358);
   U2004 : INV_X1 port map( A => n2358, ZN => n2736);
   U2005 : MUX2_X1 port map( A => n4432, B => n1706, S => n307, Z => n2359);
   U2006 : INV_X1 port map( A => n2359, ZN => n2737);
   U2007 : MUX2_X1 port map( A => n4434, B => n1741, S => n307, Z => n2360);
   U2008 : INV_X1 port map( A => n2360, ZN => n2738);
   U2009 : MUX2_X1 port map( A => n4436, B => n1777, S => n307, Z => n2361);
   U2010 : INV_X1 port map( A => n2361, ZN => n2739);
   U2011 : MUX2_X1 port map( A => n4438, B => n1813, S => n307, Z => n2362);
   U2012 : INV_X1 port map( A => n2362, ZN => n2740);
   U2013 : MUX2_X1 port map( A => n4440, B => n1849, S => n307, Z => n2363);
   U2014 : INV_X1 port map( A => n2363, ZN => n2741);
   U2015 : MUX2_X1 port map( A => n4442, B => n1885, S => n307, Z => n2364);
   U2016 : INV_X1 port map( A => n2364, ZN => n2742);
   U2017 : MUX2_X1 port map( A => n4444, B => n1921, S => n308, Z => n2365);
   U2018 : INV_X1 port map( A => n2365, ZN => n2743);
   U2019 : MUX2_X1 port map( A => n4446, B => n1957, S => n308, Z => n2366);
   U2020 : INV_X1 port map( A => n2366, ZN => n2744);
   U2021 : MUX2_X1 port map( A => n4448, B => n1992, S => n308, Z => n2367);
   U2022 : INV_X1 port map( A => n2367, ZN => n2745);
   U2023 : MUX2_X1 port map( A => n4450, B => n2027, S => n308, Z => n2368);
   U2024 : INV_X1 port map( A => n2368, ZN => n2746);
   U2025 : MUX2_X1 port map( A => n4452, B => n2063, S => n308, Z => n2369);
   U2026 : INV_X1 port map( A => n2369, ZN => n2747);
   U2027 : MUX2_X1 port map( A => n4454, B => n2099, S => n308, Z => n2370);
   U2028 : INV_X1 port map( A => n2370, ZN => n2748);
   U2029 : MUX2_X1 port map( A => n4456, B => n2135, S => n308, Z => n2371);
   U2030 : INV_X1 port map( A => n2371, ZN => n2749);
   U2031 : MUX2_X1 port map( A => n4459, B => n2182, S => n308, Z => n2373);
   U2032 : INV_X1 port map( A => n2373, ZN => n2750);
   U2033 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n2444, A3 => n2442, ZN => 
                           n4291);
   U2034 : OAI21_X1 port map( B1 => n4291, B2 => n2445, A => n84, ZN => n2374);
   U2035 : INV_X1 port map( A => n2374, ZN => n2406);
   U2036 : MUX2_X1 port map( A => n4396, B => n1062, S => n309, Z => n2375);
   U2037 : INV_X1 port map( A => n2375, ZN => n2751);
   U2038 : MUX2_X1 port map( A => n4398, B => n1100, S => n309, Z => n2376);
   U2039 : INV_X1 port map( A => n2376, ZN => n2752);
   U2040 : MUX2_X1 port map( A => n4400, B => n1136, S => n309, Z => n2377);
   U2041 : INV_X1 port map( A => n2377, ZN => n2753);
   U2042 : MUX2_X1 port map( A => n4402, B => n1172, S => n309, Z => n2378);
   U2043 : INV_X1 port map( A => n2378, ZN => n2754);
   U2044 : MUX2_X1 port map( A => n4404, B => n1208, S => n309, Z => n2379);
   U2045 : INV_X1 port map( A => n2379, ZN => n2755);
   U2046 : MUX2_X1 port map( A => n4406, B => n1244, S => n309, Z => n2380);
   U2047 : INV_X1 port map( A => n2380, ZN => n2756);
   U2048 : MUX2_X1 port map( A => n4408, B => n1280, S => n309, Z => n2381);
   U2049 : INV_X1 port map( A => n2381, ZN => n2757);
   U2050 : MUX2_X1 port map( A => n4410, B => n1316, S => n309, Z => n2382);
   U2051 : INV_X1 port map( A => n2382, ZN => n2758);
   U2052 : MUX2_X1 port map( A => n4412, B => n1352, S => n309, Z => n2383);
   U2053 : INV_X1 port map( A => n2383, ZN => n2759);
   U2054 : MUX2_X1 port map( A => n4414, B => n1387, S => n309, Z => n2384);
   U2055 : INV_X1 port map( A => n2384, ZN => n2760);
   U2056 : MUX2_X1 port map( A => n4416, B => n1422, S => n309, Z => n2385);
   U2057 : INV_X1 port map( A => n2385, ZN => n2761);
   U2058 : MUX2_X1 port map( A => n4418, B => n1457, S => n309, Z => n2386);
   U2059 : INV_X1 port map( A => n2386, ZN => n2762);
   U2060 : MUX2_X1 port map( A => n4420, B => n1492, S => n310, Z => n2387);
   U2061 : INV_X1 port map( A => n2387, ZN => n2763);
   U2062 : MUX2_X1 port map( A => n4422, B => n1527, S => n310, Z => n2388);
   U2063 : INV_X1 port map( A => n2388, ZN => n2764);
   U2064 : MUX2_X1 port map( A => n4424, B => n1563, S => n310, Z => n2389);
   U2065 : INV_X1 port map( A => n2389, ZN => n2765);
   U2066 : MUX2_X1 port map( A => n4426, B => n1598, S => n310, Z => n2390);
   U2067 : INV_X1 port map( A => n2390, ZN => n2766);
   U2068 : MUX2_X1 port map( A => n4428, B => n1633, S => n310, Z => n2391);
   U2069 : INV_X1 port map( A => n2391, ZN => n2767);
   U2070 : MUX2_X1 port map( A => n4430, B => n1669, S => n310, Z => n2392);
   U2071 : INV_X1 port map( A => n2392, ZN => n2768);
   U2072 : MUX2_X1 port map( A => n4432, B => n1705, S => n310, Z => n2393);
   U2073 : INV_X1 port map( A => n2393, ZN => n2769);
   U2074 : MUX2_X1 port map( A => n4434, B => n1740, S => n310, Z => n2394);
   U2075 : INV_X1 port map( A => n2394, ZN => n2770);
   U2076 : MUX2_X1 port map( A => n4436, B => n1776, S => n310, Z => n2395);
   U2077 : INV_X1 port map( A => n2395, ZN => n2771);
   U2078 : MUX2_X1 port map( A => n4438, B => n1812, S => n310, Z => n2396);
   U2079 : INV_X1 port map( A => n2396, ZN => n2772);
   U2080 : MUX2_X1 port map( A => n4440, B => n1848, S => n310, Z => n2397);
   U2081 : INV_X1 port map( A => n2397, ZN => n2773);
   U2082 : MUX2_X1 port map( A => n4442, B => n1884, S => n310, Z => n2398);
   U2083 : INV_X1 port map( A => n2398, ZN => n2774);
   U2084 : MUX2_X1 port map( A => n4444, B => n1920, S => n311, Z => n2399);
   U2085 : INV_X1 port map( A => n2399, ZN => n2775);
   U2086 : MUX2_X1 port map( A => n4446, B => n1956, S => n311, Z => n2400);
   U2087 : INV_X1 port map( A => n2400, ZN => n2776);
   U2088 : MUX2_X1 port map( A => n4448, B => n1991, S => n311, Z => n2401);
   U2089 : INV_X1 port map( A => n2401, ZN => n2777);
   U2090 : MUX2_X1 port map( A => n4450, B => n2026, S => n311, Z => n2402);
   U2091 : INV_X1 port map( A => n2402, ZN => n2778);
   U2092 : MUX2_X1 port map( A => n4452, B => n2062, S => n311, Z => n2403);
   U2093 : INV_X1 port map( A => n2403, ZN => n2779);
   U2094 : MUX2_X1 port map( A => n4454, B => n2098, S => n311, Z => n2404);
   U2095 : INV_X1 port map( A => n2404, ZN => n2780);
   U2096 : MUX2_X1 port map( A => n4456, B => n2134, S => n311, Z => n2405);
   U2097 : INV_X1 port map( A => n2405, ZN => n2781);
   U2098 : MUX2_X1 port map( A => n4459, B => n2180, S => n311, Z => n2407);
   U2099 : INV_X1 port map( A => n2407, ZN => n2782);
   U2100 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2444, A3 => n2443, ZN => 
                           n4358);
   U2101 : OAI21_X1 port map( B1 => n4358, B2 => n2445, A => n84, ZN => n2408);
   U2102 : INV_X1 port map( A => n2408, ZN => n2440);
   U2103 : MUX2_X1 port map( A => n4294, B => n2409, S => n312, Z => n2783);
   U2104 : MUX2_X1 port map( A => n4296, B => n2410, S => n312, Z => n2784);
   U2105 : MUX2_X1 port map( A => n4298, B => n2411, S => n312, Z => n2785);
   U2106 : MUX2_X1 port map( A => n4300, B => n2412, S => n312, Z => n2786);
   U2107 : MUX2_X1 port map( A => n4302, B => n2413, S => n312, Z => n2787);
   U2108 : MUX2_X1 port map( A => n4304, B => n2414, S => n312, Z => n2788);
   U2109 : MUX2_X1 port map( A => n4306, B => n2415, S => n312, Z => n2789);
   U2110 : MUX2_X1 port map( A => n4308, B => n2416, S => n312, Z => n2790);
   U2111 : MUX2_X1 port map( A => n4310, B => n2417, S => n312, Z => n2791);
   U2112 : MUX2_X1 port map( A => n4312, B => n2418, S => n312, Z => n2792);
   U2113 : MUX2_X1 port map( A => n4314, B => n2419, S => n312, Z => n2793);
   U2114 : MUX2_X1 port map( A => n4316, B => n2420, S => n312, Z => n2794);
   U2115 : MUX2_X1 port map( A => n4318, B => n2421, S => n313, Z => n2795);
   U2116 : MUX2_X1 port map( A => n4320, B => n2422, S => n313, Z => n2796);
   U2117 : MUX2_X1 port map( A => n4322, B => n2423, S => n313, Z => n2797);
   U2118 : MUX2_X1 port map( A => n4324, B => n2424, S => n313, Z => n2798);
   U2119 : MUX2_X1 port map( A => n4326, B => n2425, S => n313, Z => n2799);
   U2120 : MUX2_X1 port map( A => n4328, B => n2426, S => n313, Z => n2800);
   U2121 : MUX2_X1 port map( A => n4330, B => n2427, S => n313, Z => n2801);
   U2122 : MUX2_X1 port map( A => n4332, B => n2428, S => n313, Z => n2802);
   U2123 : MUX2_X1 port map( A => n4334, B => n2429, S => n313, Z => n2803);
   U2124 : MUX2_X1 port map( A => n4336, B => n2430, S => n313, Z => n2804);
   U2125 : MUX2_X1 port map( A => n4338, B => n2431, S => n313, Z => n2805);
   U2126 : MUX2_X1 port map( A => n4340, B => n2432, S => n313, Z => n2806);
   U2127 : MUX2_X1 port map( A => n4342, B => n2433, S => n314, Z => n2807);
   U2128 : MUX2_X1 port map( A => n4344, B => n2434, S => n314, Z => n2808);
   U2129 : MUX2_X1 port map( A => n4346, B => n2435, S => n314, Z => n2809);
   U2130 : MUX2_X1 port map( A => n4348, B => n2436, S => n314, Z => n2810);
   U2131 : MUX2_X1 port map( A => n4350, B => n2437, S => n314, Z => n2811);
   U2132 : MUX2_X1 port map( A => n4352, B => n2438, S => n314, Z => n2812);
   U2133 : MUX2_X1 port map( A => n4354, B => n2439, S => n314, Z => n2813);
   U2134 : MUX2_X1 port map( A => n4357, B => n2441, S => n314, Z => n2814);
   U2135 : NAND3_X1 port map( A1 => n2444, A2 => n2443, A3 => n2442, ZN => 
                           n4393);
   U2136 : OAI21_X1 port map( B1 => n4393, B2 => n2445, A => n84, ZN => n2446);
   U2137 : INV_X1 port map( A => n2446, ZN => n2478);
   U2138 : MUX2_X1 port map( A => n4294, B => n2447, S => n315, Z => n2815);
   U2139 : MUX2_X1 port map( A => n4296, B => n2448, S => n315, Z => n2816);
   U2140 : MUX2_X1 port map( A => n4298, B => n2449, S => n315, Z => n2817);
   U2141 : MUX2_X1 port map( A => n4300, B => n2450, S => n315, Z => n2818);
   U2142 : MUX2_X1 port map( A => n4302, B => n2451, S => n315, Z => n2819);
   U2143 : MUX2_X1 port map( A => n4304, B => n2452, S => n315, Z => n2820);
   U2144 : MUX2_X1 port map( A => n4306, B => n2453, S => n315, Z => n2821);
   U2145 : MUX2_X1 port map( A => n4308, B => n2454, S => n315, Z => n2822);
   U2146 : MUX2_X1 port map( A => n4310, B => n2455, S => n315, Z => n2823);
   U2147 : MUX2_X1 port map( A => n4312, B => n2456, S => n315, Z => n2824);
   U2148 : MUX2_X1 port map( A => n4314, B => n2457, S => n315, Z => n2825);
   U2149 : MUX2_X1 port map( A => n4316, B => n2458, S => n315, Z => n2826);
   U2150 : MUX2_X1 port map( A => n4318, B => n2459, S => n316, Z => n2827);
   U2151 : MUX2_X1 port map( A => n4320, B => n2460, S => n316, Z => n2828);
   U2152 : MUX2_X1 port map( A => n4322, B => n2461, S => n316, Z => n2829);
   U2153 : MUX2_X1 port map( A => n4324, B => n2462, S => n316, Z => n2830);
   U2154 : MUX2_X1 port map( A => n4326, B => n2463, S => n316, Z => n2831);
   U2155 : MUX2_X1 port map( A => n4328, B => n2464, S => n316, Z => n2832);
   U2156 : MUX2_X1 port map( A => n4330, B => n2465, S => n316, Z => n2833);
   U2157 : MUX2_X1 port map( A => n4332, B => n2466, S => n316, Z => n2834);
   U2158 : MUX2_X1 port map( A => n4334, B => n2467, S => n316, Z => n2835);
   U2159 : MUX2_X1 port map( A => n4336, B => n2468, S => n316, Z => n2836);
   U2160 : MUX2_X1 port map( A => n4338, B => n2469, S => n316, Z => n2837);
   U2161 : MUX2_X1 port map( A => n4340, B => n2470, S => n316, Z => n2838);
   U2162 : MUX2_X1 port map( A => n4342, B => n2471, S => n317, Z => n2839);
   U2163 : MUX2_X1 port map( A => n4344, B => n2472, S => n317, Z => n2840);
   U2164 : MUX2_X1 port map( A => n4346, B => n2473, S => n317, Z => n2841);
   U2165 : MUX2_X1 port map( A => n4348, B => n2474, S => n317, Z => n2842);
   U2166 : MUX2_X1 port map( A => n4350, B => n2475, S => n317, Z => n2843);
   U2167 : MUX2_X1 port map( A => n4352, B => n2476, S => n317, Z => n2844);
   U2168 : MUX2_X1 port map( A => n4354, B => n2477, S => n317, Z => n2845);
   U2169 : MUX2_X1 port map( A => n4357, B => n2479, S => n317, Z => n2846);
   U2170 : INV_X1 port map( A => ADD_WR(3), ZN => n4115);
   U2171 : NAND2_X1 port map( A1 => n16, A2 => n4115, ZN => n3806);
   U2172 : OAI21_X1 port map( B1 => n4116, B2 => n3806, A => n84, ZN => n2480);
   U2173 : INV_X1 port map( A => n2480, ZN => n2512);
   U2174 : MUX2_X1 port map( A => n4294, B => n2481, S => n318, Z => n2847);
   U2175 : MUX2_X1 port map( A => n4296, B => n2482, S => n318, Z => n2848);
   U2176 : MUX2_X1 port map( A => n4298, B => n2483, S => n318, Z => n2849);
   U2177 : MUX2_X1 port map( A => n4300, B => n2484, S => n318, Z => n2850);
   U2178 : MUX2_X1 port map( A => n4302, B => n2485, S => n318, Z => n2851);
   U2179 : MUX2_X1 port map( A => n4304, B => n2486, S => n318, Z => n2852);
   U2180 : MUX2_X1 port map( A => n4306, B => n2487, S => n318, Z => n2853);
   U2181 : MUX2_X1 port map( A => n4308, B => n2488, S => n318, Z => n2854);
   U2182 : MUX2_X1 port map( A => n4310, B => n2489, S => n318, Z => n2855);
   U2183 : MUX2_X1 port map( A => n4312, B => n2490, S => n318, Z => n2856);
   U2184 : MUX2_X1 port map( A => n4314, B => n2491, S => n318, Z => n2857);
   U2185 : MUX2_X1 port map( A => n4316, B => n2492, S => n318, Z => n2858);
   U2186 : MUX2_X1 port map( A => n4318, B => n2493, S => n319, Z => n2859);
   U2187 : MUX2_X1 port map( A => n4320, B => n2494, S => n319, Z => n2860);
   U2188 : MUX2_X1 port map( A => n4322, B => n2495, S => n319, Z => n2861);
   U2189 : MUX2_X1 port map( A => n4324, B => n2496, S => n319, Z => n2862);
   U2190 : MUX2_X1 port map( A => n4326, B => n2497, S => n319, Z => n2863);
   U2191 : MUX2_X1 port map( A => n4328, B => n2498, S => n319, Z => n2864);
   U2192 : MUX2_X1 port map( A => n4330, B => n2499, S => n319, Z => n2865);
   U2193 : MUX2_X1 port map( A => n4332, B => n2500, S => n319, Z => n2866);
   U2194 : MUX2_X1 port map( A => n4334, B => n2501, S => n319, Z => n2867);
   U2195 : MUX2_X1 port map( A => n4336, B => n2502, S => n319, Z => n2868);
   U2196 : MUX2_X1 port map( A => n4338, B => n2503, S => n319, Z => n2869);
   U2197 : MUX2_X1 port map( A => n4340, B => n2504, S => n319, Z => n2870);
   U2198 : MUX2_X1 port map( A => n4342, B => n2505, S => n320, Z => n2871);
   U2199 : MUX2_X1 port map( A => n4344, B => n2506, S => n320, Z => n2872);
   U2200 : MUX2_X1 port map( A => n4346, B => n2507, S => n320, Z => n2873);
   U2201 : MUX2_X1 port map( A => n4348, B => n2508, S => n320, Z => n2874);
   U2202 : MUX2_X1 port map( A => n4350, B => n2509, S => n320, Z => n2875);
   U2203 : MUX2_X1 port map( A => n4352, B => n2510, S => n320, Z => n2876);
   U2204 : MUX2_X1 port map( A => n4354, B => n2511, S => n320, Z => n2877);
   U2205 : MUX2_X1 port map( A => n4357, B => n2513, S => n320, Z => n2878);
   U2206 : OAI21_X1 port map( B1 => n4151, B2 => n3806, A => n83, ZN => n2514);
   U2207 : INV_X1 port map( A => n2514, ZN => n3634);
   U2208 : MUX2_X1 port map( A => n4294, B => n2515, S => n321, Z => n2879);
   U2209 : MUX2_X1 port map( A => n4296, B => n2516, S => n321, Z => n2880);
   U2210 : MUX2_X1 port map( A => n4298, B => n2517, S => n321, Z => n2881);
   U2211 : MUX2_X1 port map( A => n4300, B => n2518, S => n321, Z => n2882);
   U2212 : MUX2_X1 port map( A => n4302, B => n2519, S => n321, Z => n2883);
   U2213 : MUX2_X1 port map( A => n4304, B => n2520, S => n321, Z => n2884);
   U2214 : MUX2_X1 port map( A => n4306, B => n2521, S => n321, Z => n2885);
   U2215 : MUX2_X1 port map( A => n4308, B => n2522, S => n321, Z => n2886);
   U2216 : MUX2_X1 port map( A => n4310, B => n2523, S => n321, Z => n2887);
   U2217 : MUX2_X1 port map( A => n4312, B => n2524, S => n321, Z => n2888);
   U2218 : MUX2_X1 port map( A => n4314, B => n2525, S => n321, Z => n2889);
   U2219 : MUX2_X1 port map( A => n4316, B => n2526, S => n321, Z => n2890);
   U2220 : MUX2_X1 port map( A => n4318, B => n3615, S => n322, Z => n2891);
   U2221 : MUX2_X1 port map( A => n4320, B => n3616, S => n322, Z => n2892);
   U2222 : MUX2_X1 port map( A => n4322, B => n3617, S => n322, Z => n2893);
   U2223 : MUX2_X1 port map( A => n4324, B => n3618, S => n322, Z => n2894);
   U2224 : MUX2_X1 port map( A => n4326, B => n3619, S => n322, Z => n2895);
   U2225 : MUX2_X1 port map( A => n4328, B => n3620, S => n322, Z => n2896);
   U2226 : MUX2_X1 port map( A => n4330, B => n3621, S => n322, Z => n2897);
   U2227 : MUX2_X1 port map( A => n4332, B => n3622, S => n322, Z => n2898);
   U2228 : MUX2_X1 port map( A => n4334, B => n3623, S => n322, Z => n2899);
   U2229 : MUX2_X1 port map( A => n4336, B => n3624, S => n322, Z => n2900);
   U2230 : MUX2_X1 port map( A => n4338, B => n3625, S => n322, Z => n2901);
   U2231 : MUX2_X1 port map( A => n4340, B => n3626, S => n322, Z => n2902);
   U2232 : MUX2_X1 port map( A => n4342, B => n3627, S => n323, Z => n2903);
   U2233 : MUX2_X1 port map( A => n4344, B => n3628, S => n323, Z => n2904);
   U2234 : MUX2_X1 port map( A => n4346, B => n3629, S => n323, Z => n2905);
   U2235 : MUX2_X1 port map( A => n4348, B => n3630, S => n323, Z => n2906);
   U2236 : MUX2_X1 port map( A => n4350, B => n3631, S => n323, Z => n2907);
   U2237 : MUX2_X1 port map( A => n4352, B => n3632, S => n323, Z => n2908);
   U2238 : MUX2_X1 port map( A => n4354, B => n3633, S => n323, Z => n2909);
   U2239 : MUX2_X1 port map( A => n4357, B => n3635, S => n323, Z => n2910);
   U2240 : OAI21_X1 port map( B1 => n4186, B2 => n3806, A => n83, ZN => n3636);
   U2241 : INV_X1 port map( A => n3636, ZN => n3668);
   U2242 : MUX2_X1 port map( A => n4396, B => n1068, S => n324, Z => n3637);
   U2243 : INV_X1 port map( A => n3637, ZN => n2911);
   U2244 : MUX2_X1 port map( A => n4398, B => n1104, S => n324, Z => n3638);
   U2245 : INV_X1 port map( A => n3638, ZN => n2912);
   U2246 : MUX2_X1 port map( A => n4400, B => n1140, S => n324, Z => n3639);
   U2247 : INV_X1 port map( A => n3639, ZN => n2913);
   U2248 : MUX2_X1 port map( A => n4402, B => n1176, S => n324, Z => n3640);
   U2249 : INV_X1 port map( A => n3640, ZN => n2914);
   U2250 : MUX2_X1 port map( A => n4404, B => n1212, S => n324, Z => n3641);
   U2251 : INV_X1 port map( A => n3641, ZN => n2915);
   U2252 : MUX2_X1 port map( A => n4406, B => n1248, S => n324, Z => n3642);
   U2253 : INV_X1 port map( A => n3642, ZN => n2916);
   U2254 : MUX2_X1 port map( A => n4408, B => n1284, S => n324, Z => n3643);
   U2255 : INV_X1 port map( A => n3643, ZN => n2917);
   U2256 : MUX2_X1 port map( A => n4410, B => n1320, S => n324, Z => n3644);
   U2257 : INV_X1 port map( A => n3644, ZN => n2918);
   U2258 : MUX2_X1 port map( A => n4412, B => n1356, S => n324, Z => n3645);
   U2259 : INV_X1 port map( A => n3645, ZN => n2919);
   U2260 : MUX2_X1 port map( A => n4414, B => n1391, S => n324, Z => n3646);
   U2261 : INV_X1 port map( A => n3646, ZN => n2920);
   U2262 : MUX2_X1 port map( A => n4416, B => n1426, S => n324, Z => n3647);
   U2263 : INV_X1 port map( A => n3647, ZN => n2921);
   U2264 : MUX2_X1 port map( A => n4418, B => n1461, S => n324, Z => n3648);
   U2265 : INV_X1 port map( A => n3648, ZN => n2922);
   U2266 : MUX2_X1 port map( A => n4420, B => n1496, S => n325, Z => n3649);
   U2267 : INV_X1 port map( A => n3649, ZN => n2923);
   U2268 : MUX2_X1 port map( A => n4422, B => n1531, S => n325, Z => n3650);
   U2269 : INV_X1 port map( A => n3650, ZN => n2924);
   U2270 : MUX2_X1 port map( A => n4424, B => n1567, S => n325, Z => n3651);
   U2271 : INV_X1 port map( A => n3651, ZN => n2925);
   U2272 : MUX2_X1 port map( A => n4426, B => n1602, S => n325, Z => n3652);
   U2273 : INV_X1 port map( A => n3652, ZN => n2926);
   U2274 : MUX2_X1 port map( A => n4428, B => n1637, S => n325, Z => n3653);
   U2275 : INV_X1 port map( A => n3653, ZN => n2927);
   U2276 : MUX2_X1 port map( A => n4430, B => n1673, S => n325, Z => n3654);
   U2277 : INV_X1 port map( A => n3654, ZN => n2928);
   U2278 : MUX2_X1 port map( A => n4432, B => n1709, S => n325, Z => n3655);
   U2279 : INV_X1 port map( A => n3655, ZN => n2929);
   U2280 : MUX2_X1 port map( A => n4434, B => n1744, S => n325, Z => n3656);
   U2281 : INV_X1 port map( A => n3656, ZN => n2930);
   U2282 : MUX2_X1 port map( A => n4436, B => n1780, S => n325, Z => n3657);
   U2283 : INV_X1 port map( A => n3657, ZN => n2931);
   U2284 : MUX2_X1 port map( A => n4438, B => n1816, S => n325, Z => n3658);
   U2285 : INV_X1 port map( A => n3658, ZN => n2932);
   U2286 : MUX2_X1 port map( A => n4440, B => n1852, S => n325, Z => n3659);
   U2287 : INV_X1 port map( A => n3659, ZN => n2933);
   U2288 : MUX2_X1 port map( A => n4442, B => n1888, S => n325, Z => n3660);
   U2289 : INV_X1 port map( A => n3660, ZN => n2934);
   U2290 : MUX2_X1 port map( A => n4444, B => n1924, S => n326, Z => n3661);
   U2291 : INV_X1 port map( A => n3661, ZN => n2935);
   U2292 : MUX2_X1 port map( A => n4446, B => n1960, S => n326, Z => n3662);
   U2293 : INV_X1 port map( A => n3662, ZN => n2936);
   U2294 : MUX2_X1 port map( A => n4448, B => n1995, S => n326, Z => n3663);
   U2295 : INV_X1 port map( A => n3663, ZN => n2937);
   U2296 : MUX2_X1 port map( A => n4450, B => n2030, S => n326, Z => n3664);
   U2297 : INV_X1 port map( A => n3664, ZN => n2938);
   U2298 : MUX2_X1 port map( A => n4452, B => n2066, S => n326, Z => n3665);
   U2299 : INV_X1 port map( A => n3665, ZN => n2939);
   U2300 : MUX2_X1 port map( A => n4454, B => n2102, S => n326, Z => n3666);
   U2301 : INV_X1 port map( A => n3666, ZN => n2940);
   U2302 : MUX2_X1 port map( A => n4456, B => n2138, S => n326, Z => n3667);
   U2303 : INV_X1 port map( A => n3667, ZN => n2941);
   U2304 : MUX2_X1 port map( A => n4459, B => n2187, S => n326, Z => n3669);
   U2305 : INV_X1 port map( A => n3669, ZN => n2942);
   U2306 : OAI21_X1 port map( B1 => n4221, B2 => n3806, A => n83, ZN => n3670);
   U2307 : INV_X1 port map( A => n3670, ZN => n3702);
   U2308 : MUX2_X1 port map( A => n4396, B => n1067, S => n327, Z => n3671);
   U2309 : INV_X1 port map( A => n3671, ZN => n2943);
   U2310 : MUX2_X1 port map( A => n4398, B => n1103, S => n327, Z => n3672);
   U2311 : INV_X1 port map( A => n3672, ZN => n2944);
   U2312 : MUX2_X1 port map( A => n4400, B => n1139, S => n327, Z => n3673);
   U2313 : INV_X1 port map( A => n3673, ZN => n2945);
   U2314 : MUX2_X1 port map( A => n4402, B => n1175, S => n327, Z => n3674);
   U2315 : INV_X1 port map( A => n3674, ZN => n2946);
   U2316 : MUX2_X1 port map( A => n4404, B => n1211, S => n327, Z => n3675);
   U2317 : INV_X1 port map( A => n3675, ZN => n2947);
   U2318 : MUX2_X1 port map( A => n4406, B => n1247, S => n327, Z => n3676);
   U2319 : INV_X1 port map( A => n3676, ZN => n2948);
   U2320 : MUX2_X1 port map( A => n4408, B => n1283, S => n327, Z => n3677);
   U2321 : INV_X1 port map( A => n3677, ZN => n2949);
   U2322 : MUX2_X1 port map( A => n4410, B => n1319, S => n327, Z => n3678);
   U2323 : INV_X1 port map( A => n3678, ZN => n2950);
   U2324 : MUX2_X1 port map( A => n4412, B => n1355, S => n327, Z => n3679);
   U2325 : INV_X1 port map( A => n3679, ZN => n2951);
   U2326 : MUX2_X1 port map( A => n4414, B => n1390, S => n327, Z => n3680);
   U2327 : INV_X1 port map( A => n3680, ZN => n2952);
   U2328 : MUX2_X1 port map( A => n4416, B => n1425, S => n327, Z => n3681);
   U2329 : INV_X1 port map( A => n3681, ZN => n2953);
   U2330 : MUX2_X1 port map( A => n4418, B => n1460, S => n327, Z => n3682);
   U2331 : INV_X1 port map( A => n3682, ZN => n2954);
   U2332 : MUX2_X1 port map( A => n4420, B => n1495, S => n328, Z => n3683);
   U2333 : INV_X1 port map( A => n3683, ZN => n2955);
   U2334 : MUX2_X1 port map( A => n4422, B => n1530, S => n328, Z => n3684);
   U2335 : INV_X1 port map( A => n3684, ZN => n2956);
   U2336 : MUX2_X1 port map( A => n4424, B => n1566, S => n328, Z => n3685);
   U2337 : INV_X1 port map( A => n3685, ZN => n2957);
   U2338 : MUX2_X1 port map( A => n4426, B => n1601, S => n328, Z => n3686);
   U2339 : INV_X1 port map( A => n3686, ZN => n2958);
   U2340 : MUX2_X1 port map( A => n4428, B => n1636, S => n328, Z => n3687);
   U2341 : INV_X1 port map( A => n3687, ZN => n2959);
   U2342 : MUX2_X1 port map( A => n4430, B => n1672, S => n328, Z => n3688);
   U2343 : INV_X1 port map( A => n3688, ZN => n2960);
   U2344 : MUX2_X1 port map( A => n4432, B => n1708, S => n328, Z => n3689);
   U2345 : INV_X1 port map( A => n3689, ZN => n2961);
   U2346 : MUX2_X1 port map( A => n4434, B => n1743, S => n328, Z => n3690);
   U2347 : INV_X1 port map( A => n3690, ZN => n2962);
   U2348 : MUX2_X1 port map( A => n4436, B => n1779, S => n328, Z => n3691);
   U2349 : INV_X1 port map( A => n3691, ZN => n2963);
   U2350 : MUX2_X1 port map( A => n4438, B => n1815, S => n328, Z => n3692);
   U2351 : INV_X1 port map( A => n3692, ZN => n2964);
   U2352 : MUX2_X1 port map( A => n4440, B => n1851, S => n328, Z => n3693);
   U2353 : INV_X1 port map( A => n3693, ZN => n2965);
   U2354 : MUX2_X1 port map( A => n4442, B => n1887, S => n328, Z => n3694);
   U2355 : INV_X1 port map( A => n3694, ZN => n2966);
   U2356 : MUX2_X1 port map( A => n4444, B => n1923, S => n329, Z => n3695);
   U2357 : INV_X1 port map( A => n3695, ZN => n2967);
   U2358 : MUX2_X1 port map( A => n4446, B => n1959, S => n329, Z => n3696);
   U2359 : INV_X1 port map( A => n3696, ZN => n2968);
   U2360 : MUX2_X1 port map( A => n4448, B => n1994, S => n329, Z => n3697);
   U2361 : INV_X1 port map( A => n3697, ZN => n2969);
   U2362 : MUX2_X1 port map( A => n4450, B => n2029, S => n329, Z => n3698);
   U2363 : INV_X1 port map( A => n3698, ZN => n2970);
   U2364 : MUX2_X1 port map( A => n4452, B => n2065, S => n329, Z => n3699);
   U2365 : INV_X1 port map( A => n3699, ZN => n2971);
   U2366 : MUX2_X1 port map( A => n4454, B => n2101, S => n329, Z => n3700);
   U2367 : INV_X1 port map( A => n3700, ZN => n2972);
   U2368 : MUX2_X1 port map( A => n4456, B => n2137, S => n329, Z => n3701);
   U2369 : INV_X1 port map( A => n3701, ZN => n2973);
   U2370 : MUX2_X1 port map( A => n4459, B => n2185, S => n329, Z => n3703);
   U2371 : INV_X1 port map( A => n3703, ZN => n2974);
   U2372 : OAI21_X1 port map( B1 => n4256, B2 => n3806, A => n84, ZN => n3704);
   U2373 : INV_X1 port map( A => n3704, ZN => n3736);
   U2374 : MUX2_X1 port map( A => n4294, B => n3705, S => n330, Z => n2975);
   U2375 : MUX2_X1 port map( A => n4296, B => n3706, S => n330, Z => n2976);
   U2376 : MUX2_X1 port map( A => n4298, B => n3707, S => n330, Z => n2977);
   U2377 : MUX2_X1 port map( A => n4300, B => n3708, S => n330, Z => n2978);
   U2378 : MUX2_X1 port map( A => n4302, B => n3709, S => n330, Z => n2979);
   U2379 : MUX2_X1 port map( A => n4304, B => n3710, S => n330, Z => n2980);
   U2380 : MUX2_X1 port map( A => n4306, B => n3711, S => n330, Z => n2981);
   U2381 : MUX2_X1 port map( A => n4308, B => n3712, S => n330, Z => n2982);
   U2382 : MUX2_X1 port map( A => n4310, B => n3713, S => n330, Z => n2983);
   U2383 : MUX2_X1 port map( A => n4312, B => n3714, S => n330, Z => n2984);
   U2384 : MUX2_X1 port map( A => n4314, B => n3715, S => n330, Z => n2985);
   U2385 : MUX2_X1 port map( A => n4316, B => n3716, S => n330, Z => n2986);
   U2386 : MUX2_X1 port map( A => n4318, B => n3717, S => n331, Z => n2987);
   U2387 : MUX2_X1 port map( A => n4320, B => n3718, S => n331, Z => n2988);
   U2388 : MUX2_X1 port map( A => n4322, B => n3719, S => n331, Z => n2989);
   U2389 : MUX2_X1 port map( A => n4324, B => n3720, S => n331, Z => n2990);
   U2390 : MUX2_X1 port map( A => n4326, B => n3721, S => n331, Z => n2991);
   U2391 : MUX2_X1 port map( A => n4328, B => n3722, S => n331, Z => n2992);
   U2392 : MUX2_X1 port map( A => n4330, B => n3723, S => n331, Z => n2993);
   U2393 : MUX2_X1 port map( A => n4332, B => n3724, S => n331, Z => n2994);
   U2394 : MUX2_X1 port map( A => n4334, B => n3725, S => n331, Z => n2995);
   U2395 : MUX2_X1 port map( A => n4336, B => n3726, S => n331, Z => n2996);
   U2396 : MUX2_X1 port map( A => n4338, B => n3727, S => n331, Z => n2997);
   U2397 : MUX2_X1 port map( A => n4340, B => n3728, S => n331, Z => n2998);
   U2398 : MUX2_X1 port map( A => n4342, B => n3729, S => n332, Z => n2999);
   U2399 : MUX2_X1 port map( A => n4344, B => n3730, S => n332, Z => n3000);
   U2400 : MUX2_X1 port map( A => n4346, B => n3731, S => n332, Z => n3001);
   U2401 : MUX2_X1 port map( A => n4348, B => n3732, S => n332, Z => n3002);
   U2402 : MUX2_X1 port map( A => n4350, B => n3733, S => n332, Z => n3003);
   U2403 : MUX2_X1 port map( A => n4352, B => n3734, S => n332, Z => n3004);
   U2404 : MUX2_X1 port map( A => n4354, B => n3735, S => n332, Z => n3005);
   U2405 : MUX2_X1 port map( A => n4357, B => n3737, S => n332, Z => n3006);
   U2406 : OAI21_X1 port map( B1 => n4291, B2 => n3806, A => n83, ZN => n3738);
   U2407 : INV_X1 port map( A => n3738, ZN => n3770);
   U2408 : MUX2_X1 port map( A => n4294, B => n3739, S => n333, Z => n3007);
   U2409 : MUX2_X1 port map( A => n4296, B => n3740, S => n333, Z => n3008);
   U2410 : MUX2_X1 port map( A => n4298, B => n3741, S => n333, Z => n3009);
   U2411 : MUX2_X1 port map( A => n4300, B => n3742, S => n333, Z => n3010);
   U2412 : MUX2_X1 port map( A => n4302, B => n3743, S => n333, Z => n3011);
   U2413 : MUX2_X1 port map( A => n4304, B => n3744, S => n333, Z => n3012);
   U2414 : MUX2_X1 port map( A => n4306, B => n3745, S => n333, Z => n3013);
   U2415 : MUX2_X1 port map( A => n4308, B => n3746, S => n333, Z => n3014);
   U2416 : MUX2_X1 port map( A => n4310, B => n3747, S => n333, Z => n3015);
   U2417 : MUX2_X1 port map( A => n4312, B => n3748, S => n333, Z => n3016);
   U2418 : MUX2_X1 port map( A => n4314, B => n3749, S => n333, Z => n3017);
   U2419 : MUX2_X1 port map( A => n4316, B => n3750, S => n333, Z => n3018);
   U2420 : MUX2_X1 port map( A => n4318, B => n3751, S => n334, Z => n3019);
   U2421 : MUX2_X1 port map( A => n4320, B => n3752, S => n334, Z => n3020);
   U2422 : MUX2_X1 port map( A => n4322, B => n3753, S => n334, Z => n3021);
   U2423 : MUX2_X1 port map( A => n4324, B => n3754, S => n334, Z => n3022);
   U2424 : MUX2_X1 port map( A => n4326, B => n3755, S => n334, Z => n3023);
   U2425 : MUX2_X1 port map( A => n4328, B => n3756, S => n334, Z => n3024);
   U2426 : MUX2_X1 port map( A => n4330, B => n3757, S => n334, Z => n3025);
   U2427 : MUX2_X1 port map( A => n4332, B => n3758, S => n334, Z => n3026);
   U2428 : MUX2_X1 port map( A => n4334, B => n3759, S => n334, Z => n3027);
   U2429 : MUX2_X1 port map( A => n4336, B => n3760, S => n334, Z => n3028);
   U2430 : MUX2_X1 port map( A => n4338, B => n3761, S => n334, Z => n3029);
   U2431 : MUX2_X1 port map( A => n4340, B => n3762, S => n334, Z => n3030);
   U2432 : MUX2_X1 port map( A => n4342, B => n3763, S => n335, Z => n3031);
   U2433 : MUX2_X1 port map( A => n4344, B => n3764, S => n335, Z => n3032);
   U2434 : MUX2_X1 port map( A => n4346, B => n3765, S => n335, Z => n3033);
   U2435 : MUX2_X1 port map( A => n4348, B => n3766, S => n335, Z => n3034);
   U2436 : MUX2_X1 port map( A => n4350, B => n3767, S => n335, Z => n3035);
   U2437 : MUX2_X1 port map( A => n4352, B => n3768, S => n335, Z => n3036);
   U2438 : MUX2_X1 port map( A => n4354, B => n3769, S => n335, Z => n3037);
   U2439 : MUX2_X1 port map( A => n4357, B => n3771, S => n335, Z => n3038);
   U2440 : OAI21_X1 port map( B1 => n4358, B2 => n3806, A => n84, ZN => n3772);
   U2441 : INV_X1 port map( A => n3772, ZN => n3804);
   U2442 : MUX2_X1 port map( A => n4396, B => n1071, S => n336, Z => n3773);
   U2443 : INV_X1 port map( A => n3773, ZN => n3039);
   U2444 : MUX2_X1 port map( A => n4398, B => n1107, S => n336, Z => n3774);
   U2445 : INV_X1 port map( A => n3774, ZN => n3040);
   U2446 : MUX2_X1 port map( A => n4400, B => n1143, S => n336, Z => n3775);
   U2447 : INV_X1 port map( A => n3775, ZN => n3041);
   U2448 : MUX2_X1 port map( A => n4402, B => n1179, S => n336, Z => n3776);
   U2449 : INV_X1 port map( A => n3776, ZN => n3042);
   U2450 : MUX2_X1 port map( A => n4404, B => n1215, S => n336, Z => n3777);
   U2451 : INV_X1 port map( A => n3777, ZN => n3043);
   U2452 : MUX2_X1 port map( A => n4406, B => n1251, S => n336, Z => n3778);
   U2453 : INV_X1 port map( A => n3778, ZN => n3044);
   U2454 : MUX2_X1 port map( A => n4408, B => n1287, S => n336, Z => n3779);
   U2455 : INV_X1 port map( A => n3779, ZN => n3045);
   U2456 : MUX2_X1 port map( A => n4410, B => n1323, S => n336, Z => n3780);
   U2457 : INV_X1 port map( A => n3780, ZN => n3046);
   U2458 : MUX2_X1 port map( A => n4412, B => n1359, S => n336, Z => n3781);
   U2459 : INV_X1 port map( A => n3781, ZN => n3047);
   U2460 : MUX2_X1 port map( A => n4414, B => n1394, S => n336, Z => n3782);
   U2461 : INV_X1 port map( A => n3782, ZN => n3048);
   U2462 : MUX2_X1 port map( A => n4416, B => n1429, S => n336, Z => n3783);
   U2463 : INV_X1 port map( A => n3783, ZN => n3049);
   U2464 : MUX2_X1 port map( A => n4418, B => n1464, S => n336, Z => n3784);
   U2465 : INV_X1 port map( A => n3784, ZN => n3050);
   U2466 : MUX2_X1 port map( A => n4420, B => n1499, S => n337, Z => n3785);
   U2467 : INV_X1 port map( A => n3785, ZN => n3051);
   U2468 : MUX2_X1 port map( A => n4422, B => n1534, S => n337, Z => n3786);
   U2469 : INV_X1 port map( A => n3786, ZN => n3052);
   U2470 : MUX2_X1 port map( A => n4424, B => n1570, S => n337, Z => n3787);
   U2471 : INV_X1 port map( A => n3787, ZN => n3053);
   U2472 : MUX2_X1 port map( A => n4426, B => n1605, S => n337, Z => n3788);
   U2473 : INV_X1 port map( A => n3788, ZN => n3054);
   U2474 : MUX2_X1 port map( A => n4428, B => n1640, S => n337, Z => n3789);
   U2475 : INV_X1 port map( A => n3789, ZN => n3055);
   U2476 : MUX2_X1 port map( A => n4430, B => n1676, S => n337, Z => n3790);
   U2477 : INV_X1 port map( A => n3790, ZN => n3056);
   U2478 : MUX2_X1 port map( A => n4432, B => n1712, S => n337, Z => n3791);
   U2479 : INV_X1 port map( A => n3791, ZN => n3057);
   U2480 : MUX2_X1 port map( A => n4434, B => n1747, S => n337, Z => n3792);
   U2481 : INV_X1 port map( A => n3792, ZN => n3058);
   U2482 : MUX2_X1 port map( A => n4436, B => n1783, S => n337, Z => n3793);
   U2483 : INV_X1 port map( A => n3793, ZN => n3059);
   U2484 : MUX2_X1 port map( A => n4438, B => n1819, S => n337, Z => n3794);
   U2485 : INV_X1 port map( A => n3794, ZN => n3060);
   U2486 : MUX2_X1 port map( A => n4440, B => n1855, S => n337, Z => n3795);
   U2487 : INV_X1 port map( A => n3795, ZN => n3061);
   U2488 : MUX2_X1 port map( A => n4442, B => n1891, S => n337, Z => n3796);
   U2489 : INV_X1 port map( A => n3796, ZN => n3062);
   U2490 : MUX2_X1 port map( A => n4444, B => n1927, S => n338, Z => n3797);
   U2491 : INV_X1 port map( A => n3797, ZN => n3063);
   U2492 : MUX2_X1 port map( A => n4446, B => n1963, S => n338, Z => n3798);
   U2493 : INV_X1 port map( A => n3798, ZN => n3064);
   U2494 : MUX2_X1 port map( A => n4448, B => n1998, S => n338, Z => n3799);
   U2495 : INV_X1 port map( A => n3799, ZN => n3065);
   U2496 : MUX2_X1 port map( A => n4450, B => n2033, S => n338, Z => n3800);
   U2497 : INV_X1 port map( A => n3800, ZN => n3066);
   U2498 : MUX2_X1 port map( A => n4452, B => n2069, S => n338, Z => n3801);
   U2499 : INV_X1 port map( A => n3801, ZN => n3067);
   U2500 : MUX2_X1 port map( A => n4454, B => n2105, S => n338, Z => n3802);
   U2501 : INV_X1 port map( A => n3802, ZN => n3068);
   U2502 : MUX2_X1 port map( A => n4456, B => n2141, S => n338, Z => n3803);
   U2503 : INV_X1 port map( A => n3803, ZN => n3069);
   U2504 : MUX2_X1 port map( A => n4459, B => n2192, S => n338, Z => n3805);
   U2505 : INV_X1 port map( A => n3805, ZN => n3070);
   U2506 : OAI21_X1 port map( B1 => n4393, B2 => n3806, A => n84, ZN => n3807);
   U2507 : INV_X1 port map( A => n3807, ZN => n3839);
   U2508 : MUX2_X1 port map( A => n4396, B => n1070, S => n339, Z => n3808);
   U2509 : INV_X1 port map( A => n3808, ZN => n3071);
   U2510 : MUX2_X1 port map( A => n4398, B => n1106, S => n339, Z => n3809);
   U2511 : INV_X1 port map( A => n3809, ZN => n3072);
   U2512 : MUX2_X1 port map( A => n4400, B => n1142, S => n339, Z => n3810);
   U2513 : INV_X1 port map( A => n3810, ZN => n3073);
   U2514 : MUX2_X1 port map( A => n4402, B => n1178, S => n339, Z => n3811);
   U2515 : INV_X1 port map( A => n3811, ZN => n3074);
   U2516 : MUX2_X1 port map( A => n4404, B => n1214, S => n339, Z => n3812);
   U2517 : INV_X1 port map( A => n3812, ZN => n3075);
   U2518 : MUX2_X1 port map( A => n4406, B => n1250, S => n339, Z => n3813);
   U2519 : INV_X1 port map( A => n3813, ZN => n3076);
   U2520 : MUX2_X1 port map( A => n4408, B => n1286, S => n339, Z => n3814);
   U2521 : INV_X1 port map( A => n3814, ZN => n3077);
   U2522 : MUX2_X1 port map( A => n4410, B => n1322, S => n339, Z => n3815);
   U2523 : INV_X1 port map( A => n3815, ZN => n3078);
   U2524 : MUX2_X1 port map( A => n4412, B => n1358, S => n339, Z => n3816);
   U2525 : INV_X1 port map( A => n3816, ZN => n3079);
   U2526 : MUX2_X1 port map( A => n4414, B => n1393, S => n339, Z => n3817);
   U2527 : INV_X1 port map( A => n3817, ZN => n3080);
   U2528 : MUX2_X1 port map( A => n4416, B => n1428, S => n339, Z => n3818);
   U2529 : INV_X1 port map( A => n3818, ZN => n3081);
   U2530 : MUX2_X1 port map( A => n4418, B => n1463, S => n339, Z => n3819);
   U2531 : INV_X1 port map( A => n3819, ZN => n3082);
   U2532 : MUX2_X1 port map( A => n4420, B => n1498, S => n340, Z => n3820);
   U2533 : INV_X1 port map( A => n3820, ZN => n3083);
   U2534 : MUX2_X1 port map( A => n4422, B => n1533, S => n340, Z => n3821);
   U2535 : INV_X1 port map( A => n3821, ZN => n3084);
   U2536 : MUX2_X1 port map( A => n4424, B => n1569, S => n340, Z => n3822);
   U2537 : INV_X1 port map( A => n3822, ZN => n3085);
   U2538 : MUX2_X1 port map( A => n4426, B => n1604, S => n340, Z => n3823);
   U2539 : INV_X1 port map( A => n3823, ZN => n3086);
   U2540 : MUX2_X1 port map( A => n4428, B => n1639, S => n340, Z => n3824);
   U2541 : INV_X1 port map( A => n3824, ZN => n3087);
   U2542 : MUX2_X1 port map( A => n4430, B => n1675, S => n340, Z => n3825);
   U2543 : INV_X1 port map( A => n3825, ZN => n3088);
   U2544 : MUX2_X1 port map( A => n4432, B => n1711, S => n340, Z => n3826);
   U2545 : INV_X1 port map( A => n3826, ZN => n3089);
   U2546 : MUX2_X1 port map( A => n4434, B => n1746, S => n340, Z => n3827);
   U2547 : INV_X1 port map( A => n3827, ZN => n3090);
   U2548 : MUX2_X1 port map( A => n4436, B => n1782, S => n340, Z => n3828);
   U2549 : INV_X1 port map( A => n3828, ZN => n3091);
   U2550 : MUX2_X1 port map( A => n4438, B => n1818, S => n340, Z => n3829);
   U2551 : INV_X1 port map( A => n3829, ZN => n3092);
   U2552 : MUX2_X1 port map( A => n4440, B => n1854, S => n340, Z => n3830);
   U2553 : INV_X1 port map( A => n3830, ZN => n3093);
   U2554 : MUX2_X1 port map( A => n4442, B => n1890, S => n340, Z => n3831);
   U2555 : INV_X1 port map( A => n3831, ZN => n3094);
   U2556 : MUX2_X1 port map( A => n4444, B => n1926, S => n341, Z => n3832);
   U2557 : INV_X1 port map( A => n3832, ZN => n3095);
   U2558 : MUX2_X1 port map( A => n4446, B => n1962, S => n341, Z => n3833);
   U2559 : INV_X1 port map( A => n3833, ZN => n3096);
   U2560 : MUX2_X1 port map( A => n4448, B => n1997, S => n341, Z => n3834);
   U2561 : INV_X1 port map( A => n3834, ZN => n3097);
   U2562 : MUX2_X1 port map( A => n4450, B => n2032, S => n341, Z => n3835);
   U2563 : INV_X1 port map( A => n3835, ZN => n3098);
   U2564 : MUX2_X1 port map( A => n4452, B => n2068, S => n341, Z => n3836);
   U2565 : INV_X1 port map( A => n3836, ZN => n3099);
   U2566 : MUX2_X1 port map( A => n4454, B => n2104, S => n341, Z => n3837);
   U2567 : INV_X1 port map( A => n3837, ZN => n3100);
   U2568 : MUX2_X1 port map( A => n4456, B => n2140, S => n341, Z => n3838);
   U2569 : INV_X1 port map( A => n3838, ZN => n3101);
   U2570 : MUX2_X1 port map( A => n4459, B => n2190, S => n341, Z => n3840);
   U2571 : INV_X1 port map( A => n3840, ZN => n3102);
   U2572 : INV_X1 port map( A => ADD_WR(4), ZN => n4114);
   U2573 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => WR, A3 => n4114, ZN => 
                           n4079);
   U2574 : OAI21_X1 port map( B1 => n4116, B2 => n4079, A => n84, ZN => n3841);
   U2575 : INV_X1 port map( A => n3841, ZN => n3873);
   U2576 : MUX2_X1 port map( A => n4294, B => n3842, S => n342, Z => n3103);
   U2577 : MUX2_X1 port map( A => n4296, B => n3843, S => n342, Z => n3104);
   U2578 : MUX2_X1 port map( A => n4298, B => n3844, S => n342, Z => n3105);
   U2579 : MUX2_X1 port map( A => n4300, B => n3845, S => n342, Z => n3106);
   U2580 : MUX2_X1 port map( A => n4302, B => n3846, S => n342, Z => n3107);
   U2581 : MUX2_X1 port map( A => n4304, B => n3847, S => n342, Z => n3108);
   U2582 : MUX2_X1 port map( A => n4306, B => n3848, S => n342, Z => n3109);
   U2583 : MUX2_X1 port map( A => n4308, B => n3849, S => n342, Z => n3110);
   U2584 : MUX2_X1 port map( A => n4310, B => n3850, S => n342, Z => n3111);
   U2585 : MUX2_X1 port map( A => n4312, B => n3851, S => n342, Z => n3112);
   U2586 : MUX2_X1 port map( A => n4314, B => n3852, S => n342, Z => n3113);
   U2587 : MUX2_X1 port map( A => n4316, B => n3853, S => n342, Z => n3114);
   U2588 : MUX2_X1 port map( A => n4318, B => n3854, S => n343, Z => n3115);
   U2589 : MUX2_X1 port map( A => n4320, B => n3855, S => n343, Z => n3116);
   U2590 : MUX2_X1 port map( A => n4322, B => n3856, S => n343, Z => n3117);
   U2591 : MUX2_X1 port map( A => n4324, B => n3857, S => n343, Z => n3118);
   U2592 : MUX2_X1 port map( A => n4326, B => n3858, S => n343, Z => n3119);
   U2593 : MUX2_X1 port map( A => n4328, B => n3859, S => n343, Z => n3120);
   U2594 : MUX2_X1 port map( A => n4330, B => n3860, S => n343, Z => n3121);
   U2595 : MUX2_X1 port map( A => n4332, B => n3861, S => n343, Z => n3122);
   U2596 : MUX2_X1 port map( A => n4334, B => n3862, S => n343, Z => n3123);
   U2597 : MUX2_X1 port map( A => n4336, B => n3863, S => n343, Z => n3124);
   U2598 : MUX2_X1 port map( A => n4338, B => n3864, S => n343, Z => n3125);
   U2599 : MUX2_X1 port map( A => n4340, B => n3865, S => n343, Z => n3126);
   U2600 : MUX2_X1 port map( A => n4342, B => n3866, S => n344, Z => n3127);
   U2601 : MUX2_X1 port map( A => n4344, B => n3867, S => n344, Z => n3128);
   U2602 : MUX2_X1 port map( A => n4346, B => n3868, S => n344, Z => n3129);
   U2603 : MUX2_X1 port map( A => n4348, B => n3869, S => n344, Z => n3130);
   U2604 : MUX2_X1 port map( A => n4350, B => n3870, S => n344, Z => n3131);
   U2605 : MUX2_X1 port map( A => n4352, B => n3871, S => n344, Z => n3132);
   U2606 : MUX2_X1 port map( A => n4354, B => n3872, S => n344, Z => n3133);
   U2607 : MUX2_X1 port map( A => n4357, B => n3874, S => n344, Z => n3134);
   U2608 : OAI21_X1 port map( B1 => n4151, B2 => n4079, A => n84, ZN => n3875);
   U2609 : INV_X1 port map( A => n3875, ZN => n3907);
   U2610 : MUX2_X1 port map( A => n4294, B => n3876, S => n345, Z => n3135);
   U2611 : MUX2_X1 port map( A => n4296, B => n3877, S => n345, Z => n3136);
   U2612 : MUX2_X1 port map( A => n4298, B => n3878, S => n345, Z => n3137);
   U2613 : MUX2_X1 port map( A => n4300, B => n3879, S => n345, Z => n3138);
   U2614 : MUX2_X1 port map( A => n4302, B => n3880, S => n345, Z => n3139);
   U2615 : MUX2_X1 port map( A => n4304, B => n3881, S => n345, Z => n3140);
   U2616 : MUX2_X1 port map( A => n4306, B => n3882, S => n345, Z => n3141);
   U2617 : MUX2_X1 port map( A => n4308, B => n3883, S => n345, Z => n3142);
   U2618 : MUX2_X1 port map( A => n4310, B => n3884, S => n345, Z => n3143);
   U2619 : MUX2_X1 port map( A => n4312, B => n3885, S => n345, Z => n3144);
   U2620 : MUX2_X1 port map( A => n4314, B => n3886, S => n345, Z => n3145);
   U2621 : MUX2_X1 port map( A => n4316, B => n3887, S => n345, Z => n3146);
   U2622 : MUX2_X1 port map( A => n4318, B => n3888, S => n346, Z => n3147);
   U2623 : MUX2_X1 port map( A => n4320, B => n3889, S => n346, Z => n3148);
   U2624 : MUX2_X1 port map( A => n4322, B => n3890, S => n346, Z => n3149);
   U2625 : MUX2_X1 port map( A => n4324, B => n3891, S => n346, Z => n3150);
   U2626 : MUX2_X1 port map( A => n4326, B => n3892, S => n346, Z => n3151);
   U2627 : MUX2_X1 port map( A => n4328, B => n3893, S => n346, Z => n3152);
   U2628 : MUX2_X1 port map( A => n4330, B => n3894, S => n346, Z => n3153);
   U2629 : MUX2_X1 port map( A => n4332, B => n3895, S => n346, Z => n3154);
   U2630 : MUX2_X1 port map( A => n4334, B => n3896, S => n346, Z => n3155);
   U2631 : MUX2_X1 port map( A => n4336, B => n3897, S => n346, Z => n3156);
   U2632 : MUX2_X1 port map( A => n4338, B => n3898, S => n346, Z => n3157);
   U2633 : MUX2_X1 port map( A => n4340, B => n3899, S => n346, Z => n3158);
   U2634 : MUX2_X1 port map( A => n4342, B => n3900, S => n347, Z => n3159);
   U2635 : MUX2_X1 port map( A => n4344, B => n3901, S => n347, Z => n3160);
   U2636 : MUX2_X1 port map( A => n4346, B => n3902, S => n347, Z => n3161);
   U2637 : MUX2_X1 port map( A => n4348, B => n3903, S => n347, Z => n3162);
   U2638 : MUX2_X1 port map( A => n4350, B => n3904, S => n347, Z => n3163);
   U2639 : MUX2_X1 port map( A => n4352, B => n3905, S => n347, Z => n3164);
   U2640 : MUX2_X1 port map( A => n4354, B => n3906, S => n347, Z => n3165);
   U2641 : MUX2_X1 port map( A => n4357, B => n3908, S => n347, Z => n3166);
   U2642 : OAI21_X1 port map( B1 => n4186, B2 => n4079, A => n84, ZN => n3909);
   U2643 : INV_X1 port map( A => n3909, ZN => n3941);
   U2644 : MUX2_X1 port map( A => n4396, B => n1041, S => n348, Z => n3910);
   U2645 : INV_X1 port map( A => n3910, ZN => n3167);
   U2646 : MUX2_X1 port map( A => n4398, B => n1082, S => n348, Z => n3911);
   U2647 : INV_X1 port map( A => n3911, ZN => n3168);
   U2648 : MUX2_X1 port map( A => n4400, B => n1118, S => n348, Z => n3912);
   U2649 : INV_X1 port map( A => n3912, ZN => n3169);
   U2650 : MUX2_X1 port map( A => n4402, B => n1154, S => n348, Z => n3913);
   U2651 : INV_X1 port map( A => n3913, ZN => n3170);
   U2652 : MUX2_X1 port map( A => n4404, B => n1190, S => n348, Z => n3914);
   U2653 : INV_X1 port map( A => n3914, ZN => n3171);
   U2654 : MUX2_X1 port map( A => n4406, B => n1226, S => n348, Z => n3915);
   U2655 : INV_X1 port map( A => n3915, ZN => n3172);
   U2656 : MUX2_X1 port map( A => n4408, B => n1262, S => n348, Z => n3916);
   U2657 : INV_X1 port map( A => n3916, ZN => n3173);
   U2658 : MUX2_X1 port map( A => n4410, B => n1298, S => n348, Z => n3917);
   U2659 : INV_X1 port map( A => n3917, ZN => n3174);
   U2660 : MUX2_X1 port map( A => n4412, B => n1334, S => n348, Z => n3918);
   U2661 : INV_X1 port map( A => n3918, ZN => n3175);
   U2662 : MUX2_X1 port map( A => n4414, B => n1369, S => n348, Z => n3919);
   U2663 : INV_X1 port map( A => n3919, ZN => n3176);
   U2664 : MUX2_X1 port map( A => n4416, B => n1404, S => n348, Z => n3920);
   U2665 : INV_X1 port map( A => n3920, ZN => n3177);
   U2666 : MUX2_X1 port map( A => n4418, B => n1439, S => n348, Z => n3921);
   U2667 : INV_X1 port map( A => n3921, ZN => n3178);
   U2668 : MUX2_X1 port map( A => n4420, B => n1474, S => n349, Z => n3922);
   U2669 : INV_X1 port map( A => n3922, ZN => n3179);
   U2670 : MUX2_X1 port map( A => n4422, B => n1509, S => n349, Z => n3923);
   U2671 : INV_X1 port map( A => n3923, ZN => n3180);
   U2672 : MUX2_X1 port map( A => n4424, B => n1545, S => n349, Z => n3924);
   U2673 : INV_X1 port map( A => n3924, ZN => n3181);
   U2674 : MUX2_X1 port map( A => n4426, B => n1580, S => n349, Z => n3925);
   U2675 : INV_X1 port map( A => n3925, ZN => n3182);
   U2676 : MUX2_X1 port map( A => n4428, B => n1615, S => n349, Z => n3926);
   U2677 : INV_X1 port map( A => n3926, ZN => n3183);
   U2678 : MUX2_X1 port map( A => n4430, B => n1651, S => n349, Z => n3927);
   U2679 : INV_X1 port map( A => n3927, ZN => n3184);
   U2680 : MUX2_X1 port map( A => n4432, B => n1687, S => n349, Z => n3928);
   U2681 : INV_X1 port map( A => n3928, ZN => n3185);
   U2682 : MUX2_X1 port map( A => n4434, B => n1722, S => n349, Z => n3929);
   U2683 : INV_X1 port map( A => n3929, ZN => n3186);
   U2684 : MUX2_X1 port map( A => n4436, B => n1758, S => n349, Z => n3930);
   U2685 : INV_X1 port map( A => n3930, ZN => n3187);
   U2686 : MUX2_X1 port map( A => n4438, B => n1794, S => n349, Z => n3931);
   U2687 : INV_X1 port map( A => n3931, ZN => n3188);
   U2688 : MUX2_X1 port map( A => n4440, B => n1830, S => n349, Z => n3932);
   U2689 : INV_X1 port map( A => n3932, ZN => n3189);
   U2690 : MUX2_X1 port map( A => n4442, B => n1866, S => n349, Z => n3933);
   U2691 : INV_X1 port map( A => n3933, ZN => n3190);
   U2692 : MUX2_X1 port map( A => n4444, B => n1902, S => n350, Z => n3934);
   U2693 : INV_X1 port map( A => n3934, ZN => n3191);
   U2694 : MUX2_X1 port map( A => n4446, B => n1938, S => n350, Z => n3935);
   U2695 : INV_X1 port map( A => n3935, ZN => n3192);
   U2696 : MUX2_X1 port map( A => n4448, B => n1973, S => n350, Z => n3936);
   U2697 : INV_X1 port map( A => n3936, ZN => n3193);
   U2698 : MUX2_X1 port map( A => n4450, B => n2008, S => n350, Z => n3937);
   U2699 : INV_X1 port map( A => n3937, ZN => n3194);
   U2700 : MUX2_X1 port map( A => n4452, B => n2044, S => n350, Z => n3938);
   U2701 : INV_X1 port map( A => n3938, ZN => n3195);
   U2702 : MUX2_X1 port map( A => n4454, B => n2080, S => n350, Z => n3939);
   U2703 : INV_X1 port map( A => n3939, ZN => n3196);
   U2704 : MUX2_X1 port map( A => n4456, B => n2116, S => n350, Z => n3940);
   U2705 : INV_X1 port map( A => n3940, ZN => n3197);
   U2706 : MUX2_X1 port map( A => n4459, B => n2153, S => n350, Z => n3942);
   U2707 : INV_X1 port map( A => n3942, ZN => n3198);
   U2708 : OAI21_X1 port map( B1 => n4221, B2 => n4079, A => n84, ZN => n3943);
   U2709 : INV_X1 port map( A => n3943, ZN => n3975);
   U2710 : MUX2_X1 port map( A => n4396, B => n1040, S => n351, Z => n3944);
   U2711 : INV_X1 port map( A => n3944, ZN => n3199);
   U2712 : MUX2_X1 port map( A => n4398, B => n1081, S => n351, Z => n3945);
   U2713 : INV_X1 port map( A => n3945, ZN => n3200);
   U2714 : MUX2_X1 port map( A => n4400, B => n1117, S => n351, Z => n3946);
   U2715 : INV_X1 port map( A => n3946, ZN => n3201);
   U2716 : MUX2_X1 port map( A => n4402, B => n1153, S => n351, Z => n3947);
   U2717 : INV_X1 port map( A => n3947, ZN => n3202);
   U2718 : MUX2_X1 port map( A => n4404, B => n1189, S => n351, Z => n3948);
   U2719 : INV_X1 port map( A => n3948, ZN => n3203);
   U2720 : MUX2_X1 port map( A => n4406, B => n1225, S => n351, Z => n3949);
   U2721 : INV_X1 port map( A => n3949, ZN => n3204);
   U2722 : MUX2_X1 port map( A => n4408, B => n1261, S => n351, Z => n3950);
   U2723 : INV_X1 port map( A => n3950, ZN => n3205);
   U2724 : MUX2_X1 port map( A => n4410, B => n1297, S => n351, Z => n3951);
   U2725 : INV_X1 port map( A => n3951, ZN => n3206);
   U2726 : MUX2_X1 port map( A => n4412, B => n1333, S => n351, Z => n3952);
   U2727 : INV_X1 port map( A => n3952, ZN => n3207);
   U2728 : MUX2_X1 port map( A => n4414, B => n1368, S => n351, Z => n3953);
   U2729 : INV_X1 port map( A => n3953, ZN => n3208);
   U2730 : MUX2_X1 port map( A => n4416, B => n1403, S => n351, Z => n3954);
   U2731 : INV_X1 port map( A => n3954, ZN => n3209);
   U2732 : MUX2_X1 port map( A => n4418, B => n1438, S => n351, Z => n3955);
   U2733 : INV_X1 port map( A => n3955, ZN => n3210);
   U2734 : MUX2_X1 port map( A => n4420, B => n1473, S => n352, Z => n3956);
   U2735 : INV_X1 port map( A => n3956, ZN => n3211);
   U2736 : MUX2_X1 port map( A => n4422, B => n1508, S => n352, Z => n3957);
   U2737 : INV_X1 port map( A => n3957, ZN => n3212);
   U2738 : MUX2_X1 port map( A => n4424, B => n1544, S => n352, Z => n3958);
   U2739 : INV_X1 port map( A => n3958, ZN => n3213);
   U2740 : MUX2_X1 port map( A => n4426, B => n1579, S => n352, Z => n3959);
   U2741 : INV_X1 port map( A => n3959, ZN => n3214);
   U2742 : MUX2_X1 port map( A => n4428, B => n1614, S => n352, Z => n3960);
   U2743 : INV_X1 port map( A => n3960, ZN => n3215);
   U2744 : MUX2_X1 port map( A => n4430, B => n1650, S => n352, Z => n3961);
   U2745 : INV_X1 port map( A => n3961, ZN => n3216);
   U2746 : MUX2_X1 port map( A => n4432, B => n1686, S => n352, Z => n3962);
   U2747 : INV_X1 port map( A => n3962, ZN => n3217);
   U2748 : MUX2_X1 port map( A => n4434, B => n1721, S => n352, Z => n3963);
   U2749 : INV_X1 port map( A => n3963, ZN => n3218);
   U2750 : MUX2_X1 port map( A => n4436, B => n1757, S => n352, Z => n3964);
   U2751 : INV_X1 port map( A => n3964, ZN => n3219);
   U2752 : MUX2_X1 port map( A => n4438, B => n1793, S => n352, Z => n3965);
   U2753 : INV_X1 port map( A => n3965, ZN => n3220);
   U2754 : MUX2_X1 port map( A => n4440, B => n1829, S => n352, Z => n3966);
   U2755 : INV_X1 port map( A => n3966, ZN => n3221);
   U2756 : MUX2_X1 port map( A => n4442, B => n1865, S => n352, Z => n3967);
   U2757 : INV_X1 port map( A => n3967, ZN => n3222);
   U2758 : MUX2_X1 port map( A => n4444, B => n1901, S => n353, Z => n3968);
   U2759 : INV_X1 port map( A => n3968, ZN => n3223);
   U2760 : MUX2_X1 port map( A => n4446, B => n1937, S => n353, Z => n3969);
   U2761 : INV_X1 port map( A => n3969, ZN => n3224);
   U2762 : MUX2_X1 port map( A => n4448, B => n1972, S => n353, Z => n3970);
   U2763 : INV_X1 port map( A => n3970, ZN => n3225);
   U2764 : MUX2_X1 port map( A => n4450, B => n2007, S => n353, Z => n3971);
   U2765 : INV_X1 port map( A => n3971, ZN => n3226);
   U2766 : MUX2_X1 port map( A => n4452, B => n2043, S => n353, Z => n3972);
   U2767 : INV_X1 port map( A => n3972, ZN => n3227);
   U2768 : MUX2_X1 port map( A => n4454, B => n2079, S => n353, Z => n3973);
   U2769 : INV_X1 port map( A => n3973, ZN => n3228);
   U2770 : MUX2_X1 port map( A => n4456, B => n2115, S => n353, Z => n3974);
   U2771 : INV_X1 port map( A => n3974, ZN => n3229);
   U2772 : MUX2_X1 port map( A => n4459, B => n2151, S => n353, Z => n3976);
   U2773 : INV_X1 port map( A => n3976, ZN => n3230);
   U2774 : OAI21_X1 port map( B1 => n4256, B2 => n4079, A => n83, ZN => n3977);
   U2775 : INV_X1 port map( A => n3977, ZN => n4009);
   U2776 : MUX2_X1 port map( A => n4294, B => n3978, S => n354, Z => n3231);
   U2777 : MUX2_X1 port map( A => n4296, B => n3979, S => n354, Z => n3232);
   U2778 : MUX2_X1 port map( A => n4298, B => n3980, S => n354, Z => n3233);
   U2779 : MUX2_X1 port map( A => n4300, B => n3981, S => n354, Z => n3234);
   U2780 : MUX2_X1 port map( A => n4302, B => n3982, S => n354, Z => n3235);
   U2781 : MUX2_X1 port map( A => n4304, B => n3983, S => n354, Z => n3236);
   U2782 : MUX2_X1 port map( A => n4306, B => n3984, S => n354, Z => n3237);
   U2783 : MUX2_X1 port map( A => n4308, B => n3985, S => n354, Z => n3238);
   U2784 : MUX2_X1 port map( A => n4310, B => n3986, S => n354, Z => n3239);
   U2785 : MUX2_X1 port map( A => n4312, B => n3987, S => n354, Z => n3240);
   U2786 : MUX2_X1 port map( A => n4314, B => n3988, S => n354, Z => n3241);
   U2787 : MUX2_X1 port map( A => n4316, B => n3989, S => n354, Z => n3242);
   U2788 : MUX2_X1 port map( A => n4318, B => n3990, S => n355, Z => n3243);
   U2789 : MUX2_X1 port map( A => n4320, B => n3991, S => n355, Z => n3244);
   U2790 : MUX2_X1 port map( A => n4322, B => n3992, S => n355, Z => n3245);
   U2791 : MUX2_X1 port map( A => n4324, B => n3993, S => n355, Z => n3246);
   U2792 : MUX2_X1 port map( A => n4326, B => n3994, S => n355, Z => n3247);
   U2793 : MUX2_X1 port map( A => n4328, B => n3995, S => n355, Z => n3248);
   U2794 : MUX2_X1 port map( A => n4330, B => n3996, S => n355, Z => n3249);
   U2795 : MUX2_X1 port map( A => n4332, B => n3997, S => n355, Z => n3250);
   U2796 : MUX2_X1 port map( A => n4334, B => n3998, S => n355, Z => n3251);
   U2797 : MUX2_X1 port map( A => n4336, B => n3999, S => n355, Z => n3252);
   U2798 : MUX2_X1 port map( A => n4338, B => n4000, S => n355, Z => n3253);
   U2799 : MUX2_X1 port map( A => n4340, B => n4001, S => n355, Z => n3254);
   U2800 : MUX2_X1 port map( A => n4342, B => n4002, S => n356, Z => n3255);
   U2801 : MUX2_X1 port map( A => n4344, B => n4003, S => n356, Z => n3256);
   U2802 : MUX2_X1 port map( A => n4346, B => n4004, S => n356, Z => n3257);
   U2803 : MUX2_X1 port map( A => n4348, B => n4005, S => n356, Z => n3258);
   U2804 : MUX2_X1 port map( A => n4350, B => n4006, S => n356, Z => n3259);
   U2805 : MUX2_X1 port map( A => n4352, B => n4007, S => n356, Z => n3260);
   U2806 : MUX2_X1 port map( A => n4354, B => n4008, S => n356, Z => n3261);
   U2807 : MUX2_X1 port map( A => n4357, B => n4010, S => n356, Z => n3262);
   U2808 : OAI21_X1 port map( B1 => n4291, B2 => n4079, A => n83, ZN => n4011);
   U2809 : INV_X1 port map( A => n4011, ZN => n4043);
   U2810 : MUX2_X1 port map( A => n4294, B => n4012, S => n357, Z => n3263);
   U2811 : MUX2_X1 port map( A => n4296, B => n4013, S => n357, Z => n3264);
   U2812 : MUX2_X1 port map( A => n4298, B => n4014, S => n357, Z => n3265);
   U2813 : MUX2_X1 port map( A => n4300, B => n4015, S => n357, Z => n3266);
   U2814 : MUX2_X1 port map( A => n4302, B => n4016, S => n357, Z => n3267);
   U2815 : MUX2_X1 port map( A => n4304, B => n4017, S => n357, Z => n3268);
   U2816 : MUX2_X1 port map( A => n4306, B => n4018, S => n357, Z => n3269);
   U2817 : MUX2_X1 port map( A => n4308, B => n4019, S => n357, Z => n3270);
   U2818 : MUX2_X1 port map( A => n4310, B => n4020, S => n357, Z => n3271);
   U2819 : MUX2_X1 port map( A => n4312, B => n4021, S => n357, Z => n3272);
   U2820 : MUX2_X1 port map( A => n4314, B => n4022, S => n357, Z => n3273);
   U2821 : MUX2_X1 port map( A => n4316, B => n4023, S => n357, Z => n3274);
   U2822 : MUX2_X1 port map( A => n4318, B => n4024, S => n358, Z => n3275);
   U2823 : MUX2_X1 port map( A => n4320, B => n4025, S => n358, Z => n3276);
   U2824 : MUX2_X1 port map( A => n4322, B => n4026, S => n358, Z => n3277);
   U2825 : MUX2_X1 port map( A => n4324, B => n4027, S => n358, Z => n3278);
   U2826 : MUX2_X1 port map( A => n4326, B => n4028, S => n358, Z => n3279);
   U2827 : MUX2_X1 port map( A => n4328, B => n4029, S => n358, Z => n3280);
   U2828 : MUX2_X1 port map( A => n4330, B => n4030, S => n358, Z => n3281);
   U2829 : MUX2_X1 port map( A => n4332, B => n4031, S => n358, Z => n3282);
   U2830 : MUX2_X1 port map( A => n4334, B => n4032, S => n358, Z => n3283);
   U2831 : MUX2_X1 port map( A => n4336, B => n4033, S => n358, Z => n3284);
   U2832 : MUX2_X1 port map( A => n4338, B => n4034, S => n358, Z => n3285);
   U2833 : MUX2_X1 port map( A => n4340, B => n4035, S => n358, Z => n3286);
   U2834 : MUX2_X1 port map( A => n4342, B => n4036, S => n359, Z => n3287);
   U2835 : MUX2_X1 port map( A => n4344, B => n4037, S => n359, Z => n3288);
   U2836 : MUX2_X1 port map( A => n4346, B => n4038, S => n359, Z => n3289);
   U2837 : MUX2_X1 port map( A => n4348, B => n4039, S => n359, Z => n3290);
   U2838 : MUX2_X1 port map( A => n4350, B => n4040, S => n359, Z => n3291);
   U2839 : MUX2_X1 port map( A => n4352, B => n4041, S => n359, Z => n3292);
   U2840 : MUX2_X1 port map( A => n4354, B => n4042, S => n359, Z => n3293);
   U2841 : MUX2_X1 port map( A => n4357, B => n4044, S => n359, Z => n3294);
   U2842 : OAI21_X1 port map( B1 => n4358, B2 => n4079, A => n83, ZN => n4045);
   U2843 : INV_X1 port map( A => n4045, ZN => n4077);
   U2844 : MUX2_X1 port map( A => n4396, B => n1046, S => n360, Z => n4046);
   U2845 : INV_X1 port map( A => n4046, ZN => n3295);
   U2846 : MUX2_X1 port map( A => n4398, B => n1085, S => n360, Z => n4047);
   U2847 : INV_X1 port map( A => n4047, ZN => n3296);
   U2848 : MUX2_X1 port map( A => n4400, B => n1121, S => n360, Z => n4048);
   U2849 : INV_X1 port map( A => n4048, ZN => n3297);
   U2850 : MUX2_X1 port map( A => n4402, B => n1157, S => n360, Z => n4049);
   U2851 : INV_X1 port map( A => n4049, ZN => n3298);
   U2852 : MUX2_X1 port map( A => n4404, B => n1193, S => n360, Z => n4050);
   U2853 : INV_X1 port map( A => n4050, ZN => n3299);
   U2854 : MUX2_X1 port map( A => n4406, B => n1229, S => n360, Z => n4051);
   U2855 : INV_X1 port map( A => n4051, ZN => n3300);
   U2856 : MUX2_X1 port map( A => n4408, B => n1265, S => n360, Z => n4052);
   U2857 : INV_X1 port map( A => n4052, ZN => n3301);
   U2858 : MUX2_X1 port map( A => n4410, B => n1301, S => n360, Z => n4053);
   U2859 : INV_X1 port map( A => n4053, ZN => n3302);
   U2860 : MUX2_X1 port map( A => n4412, B => n1337, S => n360, Z => n4054);
   U2861 : INV_X1 port map( A => n4054, ZN => n3303);
   U2862 : MUX2_X1 port map( A => n4414, B => n1372, S => n360, Z => n4055);
   U2863 : INV_X1 port map( A => n4055, ZN => n3304);
   U2864 : MUX2_X1 port map( A => n4416, B => n1407, S => n360, Z => n4056);
   U2865 : INV_X1 port map( A => n4056, ZN => n3305);
   U2866 : MUX2_X1 port map( A => n4418, B => n1442, S => n360, Z => n4057);
   U2867 : INV_X1 port map( A => n4057, ZN => n3306);
   U2868 : MUX2_X1 port map( A => n4420, B => n1477, S => n361, Z => n4058);
   U2869 : INV_X1 port map( A => n4058, ZN => n3307);
   U2870 : MUX2_X1 port map( A => n4422, B => n1512, S => n361, Z => n4059);
   U2871 : INV_X1 port map( A => n4059, ZN => n3308);
   U2872 : MUX2_X1 port map( A => n4424, B => n1548, S => n361, Z => n4060);
   U2873 : INV_X1 port map( A => n4060, ZN => n3309);
   U2874 : MUX2_X1 port map( A => n4426, B => n1583, S => n361, Z => n4061);
   U2875 : INV_X1 port map( A => n4061, ZN => n3310);
   U2876 : MUX2_X1 port map( A => n4428, B => n1618, S => n361, Z => n4062);
   U2877 : INV_X1 port map( A => n4062, ZN => n3311);
   U2878 : MUX2_X1 port map( A => n4430, B => n1654, S => n361, Z => n4063);
   U2879 : INV_X1 port map( A => n4063, ZN => n3312);
   U2880 : MUX2_X1 port map( A => n4432, B => n1690, S => n361, Z => n4064);
   U2881 : INV_X1 port map( A => n4064, ZN => n3313);
   U2882 : MUX2_X1 port map( A => n4434, B => n1725, S => n361, Z => n4065);
   U2883 : INV_X1 port map( A => n4065, ZN => n3314);
   U2884 : MUX2_X1 port map( A => n4436, B => n1761, S => n361, Z => n4066);
   U2885 : INV_X1 port map( A => n4066, ZN => n3315);
   U2886 : MUX2_X1 port map( A => n4438, B => n1797, S => n361, Z => n4067);
   U2887 : INV_X1 port map( A => n4067, ZN => n3316);
   U2888 : MUX2_X1 port map( A => n4440, B => n1833, S => n361, Z => n4068);
   U2889 : INV_X1 port map( A => n4068, ZN => n3317);
   U2890 : MUX2_X1 port map( A => n4442, B => n1869, S => n361, Z => n4069);
   U2891 : INV_X1 port map( A => n4069, ZN => n3318);
   U2892 : MUX2_X1 port map( A => n4444, B => n1905, S => n362, Z => n4070);
   U2893 : INV_X1 port map( A => n4070, ZN => n3319);
   U2894 : MUX2_X1 port map( A => n4446, B => n1941, S => n362, Z => n4071);
   U2895 : INV_X1 port map( A => n4071, ZN => n3320);
   U2896 : MUX2_X1 port map( A => n4448, B => n1976, S => n362, Z => n4072);
   U2897 : INV_X1 port map( A => n4072, ZN => n3321);
   U2898 : MUX2_X1 port map( A => n4450, B => n2011, S => n362, Z => n4073);
   U2899 : INV_X1 port map( A => n4073, ZN => n3322);
   U2900 : MUX2_X1 port map( A => n4452, B => n2047, S => n362, Z => n4074);
   U2901 : INV_X1 port map( A => n4074, ZN => n3323);
   U2902 : MUX2_X1 port map( A => n4454, B => n2083, S => n362, Z => n4075);
   U2903 : INV_X1 port map( A => n4075, ZN => n3324);
   U2904 : MUX2_X1 port map( A => n4456, B => n2119, S => n362, Z => n4076);
   U2905 : INV_X1 port map( A => n4076, ZN => n3325);
   U2906 : MUX2_X1 port map( A => n4459, B => n2158, S => n362, Z => n4078);
   U2907 : INV_X1 port map( A => n4078, ZN => n3326);
   U2908 : OAI21_X1 port map( B1 => n4393, B2 => n4079, A => n83, ZN => n4080);
   U2909 : INV_X1 port map( A => n4080, ZN => n4112);
   U2910 : MUX2_X1 port map( A => n4396, B => n1045, S => n363, Z => n4081);
   U2911 : INV_X1 port map( A => n4081, ZN => n3327);
   U2912 : MUX2_X1 port map( A => n4398, B => n1084, S => n363, Z => n4082);
   U2913 : INV_X1 port map( A => n4082, ZN => n3328);
   U2914 : MUX2_X1 port map( A => n4400, B => n1120, S => n363, Z => n4083);
   U2915 : INV_X1 port map( A => n4083, ZN => n3329);
   U2916 : MUX2_X1 port map( A => n4402, B => n1156, S => n363, Z => n4084);
   U2917 : INV_X1 port map( A => n4084, ZN => n3330);
   U2918 : MUX2_X1 port map( A => n4404, B => n1192, S => n363, Z => n4085);
   U2919 : INV_X1 port map( A => n4085, ZN => n3331);
   U2920 : MUX2_X1 port map( A => n4406, B => n1228, S => n363, Z => n4086);
   U2921 : INV_X1 port map( A => n4086, ZN => n3332);
   U2922 : MUX2_X1 port map( A => n4408, B => n1264, S => n363, Z => n4087);
   U2923 : INV_X1 port map( A => n4087, ZN => n3333);
   U2924 : MUX2_X1 port map( A => n4410, B => n1300, S => n363, Z => n4088);
   U2925 : INV_X1 port map( A => n4088, ZN => n3334);
   U2926 : MUX2_X1 port map( A => n4412, B => n1336, S => n363, Z => n4089);
   U2927 : INV_X1 port map( A => n4089, ZN => n3335);
   U2928 : MUX2_X1 port map( A => n4414, B => n1371, S => n363, Z => n4090);
   U2929 : INV_X1 port map( A => n4090, ZN => n3336);
   U2930 : MUX2_X1 port map( A => n4416, B => n1406, S => n363, Z => n4091);
   U2931 : INV_X1 port map( A => n4091, ZN => n3337);
   U2932 : MUX2_X1 port map( A => n4418, B => n1441, S => n363, Z => n4092);
   U2933 : INV_X1 port map( A => n4092, ZN => n3338);
   U2934 : MUX2_X1 port map( A => n4420, B => n1476, S => n364, Z => n4093);
   U2935 : INV_X1 port map( A => n4093, ZN => n3339);
   U2936 : MUX2_X1 port map( A => n4422, B => n1511, S => n364, Z => n4094);
   U2937 : INV_X1 port map( A => n4094, ZN => n3340);
   U2938 : MUX2_X1 port map( A => n4424, B => n1547, S => n364, Z => n4095);
   U2939 : INV_X1 port map( A => n4095, ZN => n3341);
   U2940 : MUX2_X1 port map( A => n4426, B => n1582, S => n364, Z => n4096);
   U2941 : INV_X1 port map( A => n4096, ZN => n3342);
   U2942 : MUX2_X1 port map( A => n4428, B => n1617, S => n364, Z => n4097);
   U2943 : INV_X1 port map( A => n4097, ZN => n3343);
   U2944 : MUX2_X1 port map( A => n4430, B => n1653, S => n364, Z => n4098);
   U2945 : INV_X1 port map( A => n4098, ZN => n3344);
   U2946 : MUX2_X1 port map( A => n4432, B => n1689, S => n364, Z => n4099);
   U2947 : INV_X1 port map( A => n4099, ZN => n3345);
   U2948 : MUX2_X1 port map( A => n4434, B => n1724, S => n364, Z => n4100);
   U2949 : INV_X1 port map( A => n4100, ZN => n3346);
   U2950 : MUX2_X1 port map( A => n4436, B => n1760, S => n364, Z => n4101);
   U2951 : INV_X1 port map( A => n4101, ZN => n3347);
   U2952 : MUX2_X1 port map( A => n4438, B => n1796, S => n364, Z => n4102);
   U2953 : INV_X1 port map( A => n4102, ZN => n3348);
   U2954 : MUX2_X1 port map( A => n4440, B => n1832, S => n364, Z => n4103);
   U2955 : INV_X1 port map( A => n4103, ZN => n3349);
   U2956 : MUX2_X1 port map( A => n4442, B => n1868, S => n364, Z => n4104);
   U2957 : INV_X1 port map( A => n4104, ZN => n3350);
   U2958 : MUX2_X1 port map( A => n4444, B => n1904, S => n365, Z => n4105);
   U2959 : INV_X1 port map( A => n4105, ZN => n3351);
   U2960 : MUX2_X1 port map( A => n4446, B => n1940, S => n365, Z => n4106);
   U2961 : INV_X1 port map( A => n4106, ZN => n3352);
   U2962 : MUX2_X1 port map( A => n4448, B => n1975, S => n365, Z => n4107);
   U2963 : INV_X1 port map( A => n4107, ZN => n3353);
   U2964 : MUX2_X1 port map( A => n4450, B => n2010, S => n365, Z => n4108);
   U2965 : INV_X1 port map( A => n4108, ZN => n3354);
   U2966 : MUX2_X1 port map( A => n4452, B => n2046, S => n365, Z => n4109);
   U2967 : INV_X1 port map( A => n4109, ZN => n3355);
   U2968 : MUX2_X1 port map( A => n4454, B => n2082, S => n365, Z => n4110);
   U2969 : INV_X1 port map( A => n4110, ZN => n3356);
   U2970 : MUX2_X1 port map( A => n4456, B => n2118, S => n365, Z => n4111);
   U2971 : INV_X1 port map( A => n4111, ZN => n3357);
   U2972 : MUX2_X1 port map( A => n4459, B => n2156, S => n365, Z => n4113);
   U2973 : INV_X1 port map( A => n4113, ZN => n3358);
   U2974 : NAND3_X1 port map( A1 => WR, A2 => n4115, A3 => n4114, ZN => n4394);
   U2975 : OAI21_X1 port map( B1 => n4394, B2 => n4116, A => n83, ZN => n4117);
   U2976 : INV_X1 port map( A => n4117, ZN => n4149);
   U2977 : MUX2_X1 port map( A => n4294, B => n4118, S => n366, Z => n3359);
   U2978 : MUX2_X1 port map( A => n4296, B => n4119, S => n366, Z => n3360);
   U2979 : MUX2_X1 port map( A => n4298, B => n4120, S => n366, Z => n3361);
   U2980 : MUX2_X1 port map( A => n4300, B => n4121, S => n366, Z => n3362);
   U2981 : MUX2_X1 port map( A => n4302, B => n4122, S => n366, Z => n3363);
   U2982 : MUX2_X1 port map( A => n4304, B => n4123, S => n366, Z => n3364);
   U2983 : MUX2_X1 port map( A => n4306, B => n4124, S => n366, Z => n3365);
   U2984 : MUX2_X1 port map( A => n4308, B => n4125, S => n366, Z => n3366);
   U2985 : MUX2_X1 port map( A => n4310, B => n4126, S => n366, Z => n3367);
   U2986 : MUX2_X1 port map( A => n4312, B => n4127, S => n366, Z => n3368);
   U2987 : MUX2_X1 port map( A => n4314, B => n4128, S => n366, Z => n3369);
   U2988 : MUX2_X1 port map( A => n4316, B => n4129, S => n366, Z => n3370);
   U2989 : MUX2_X1 port map( A => n4318, B => n4130, S => n367, Z => n3371);
   U2990 : MUX2_X1 port map( A => n4320, B => n4131, S => n367, Z => n3372);
   U2991 : MUX2_X1 port map( A => n4322, B => n4132, S => n367, Z => n3373);
   U2992 : MUX2_X1 port map( A => n4324, B => n4133, S => n367, Z => n3374);
   U2993 : MUX2_X1 port map( A => n4326, B => n4134, S => n367, Z => n3375);
   U2994 : MUX2_X1 port map( A => n4328, B => n4135, S => n367, Z => n3376);
   U2995 : MUX2_X1 port map( A => n4330, B => n4136, S => n367, Z => n3377);
   U2996 : MUX2_X1 port map( A => n4332, B => n4137, S => n367, Z => n3378);
   U2997 : MUX2_X1 port map( A => n4334, B => n4138, S => n367, Z => n3379);
   U2998 : MUX2_X1 port map( A => n4336, B => n4139, S => n367, Z => n3380);
   U2999 : MUX2_X1 port map( A => n4338, B => n4140, S => n367, Z => n3381);
   U3000 : MUX2_X1 port map( A => n4340, B => n4141, S => n367, Z => n3382);
   U3001 : MUX2_X1 port map( A => n4342, B => n4142, S => n368, Z => n3383);
   U3002 : MUX2_X1 port map( A => n4344, B => n4143, S => n368, Z => n3384);
   U3003 : MUX2_X1 port map( A => n4346, B => n4144, S => n368, Z => n3385);
   U3004 : MUX2_X1 port map( A => n4348, B => n4145, S => n368, Z => n3386);
   U3005 : MUX2_X1 port map( A => n4350, B => n4146, S => n368, Z => n3387);
   U3006 : MUX2_X1 port map( A => n4352, B => n4147, S => n368, Z => n3388);
   U3007 : MUX2_X1 port map( A => n4354, B => n4148, S => n368, Z => n3389);
   U3008 : MUX2_X1 port map( A => n4357, B => n4150, S => n368, Z => n3390);
   U3009 : OAI21_X1 port map( B1 => n4394, B2 => n4151, A => n84, ZN => n4152);
   U3010 : INV_X1 port map( A => n4152, ZN => n4184);
   U3011 : MUX2_X1 port map( A => n4294, B => n4153, S => n369, Z => n3391);
   U3012 : MUX2_X1 port map( A => n4296, B => n4154, S => n369, Z => n3392);
   U3013 : MUX2_X1 port map( A => n4298, B => n4155, S => n369, Z => n3393);
   U3014 : MUX2_X1 port map( A => n4300, B => n4156, S => n369, Z => n3394);
   U3015 : MUX2_X1 port map( A => n4302, B => n4157, S => n369, Z => n3395);
   U3016 : MUX2_X1 port map( A => n4304, B => n4158, S => n369, Z => n3396);
   U3017 : MUX2_X1 port map( A => n4306, B => n4159, S => n369, Z => n3397);
   U3018 : MUX2_X1 port map( A => n4308, B => n4160, S => n369, Z => n3398);
   U3019 : MUX2_X1 port map( A => n4310, B => n4161, S => n369, Z => n3399);
   U3020 : MUX2_X1 port map( A => n4312, B => n4162, S => n369, Z => n3400);
   U3021 : MUX2_X1 port map( A => n4314, B => n4163, S => n369, Z => n3401);
   U3022 : MUX2_X1 port map( A => n4316, B => n4164, S => n369, Z => n3402);
   U3023 : MUX2_X1 port map( A => n4318, B => n4165, S => n370, Z => n3403);
   U3024 : MUX2_X1 port map( A => n4320, B => n4166, S => n370, Z => n3404);
   U3025 : MUX2_X1 port map( A => n4322, B => n4167, S => n370, Z => n3405);
   U3026 : MUX2_X1 port map( A => n4324, B => n4168, S => n370, Z => n3406);
   U3027 : MUX2_X1 port map( A => n4326, B => n4169, S => n370, Z => n3407);
   U3028 : MUX2_X1 port map( A => n4328, B => n4170, S => n370, Z => n3408);
   U3029 : MUX2_X1 port map( A => n4330, B => n4171, S => n370, Z => n3409);
   U3030 : MUX2_X1 port map( A => n4332, B => n4172, S => n370, Z => n3410);
   U3031 : MUX2_X1 port map( A => n4334, B => n4173, S => n370, Z => n3411);
   U3032 : MUX2_X1 port map( A => n4336, B => n4174, S => n370, Z => n3412);
   U3033 : MUX2_X1 port map( A => n4338, B => n4175, S => n370, Z => n3413);
   U3034 : MUX2_X1 port map( A => n4340, B => n4176, S => n370, Z => n3414);
   U3035 : MUX2_X1 port map( A => n4342, B => n4177, S => n371, Z => n3415);
   U3036 : MUX2_X1 port map( A => n4344, B => n4178, S => n371, Z => n3416);
   U3037 : MUX2_X1 port map( A => n4346, B => n4179, S => n371, Z => n3417);
   U3038 : MUX2_X1 port map( A => n4348, B => n4180, S => n371, Z => n3418);
   U3039 : MUX2_X1 port map( A => n4350, B => n4181, S => n371, Z => n3419);
   U3040 : MUX2_X1 port map( A => n4352, B => n4182, S => n371, Z => n3420);
   U3041 : MUX2_X1 port map( A => n4354, B => n4183, S => n371, Z => n3421);
   U3042 : MUX2_X1 port map( A => n4357, B => n4185, S => n371, Z => n3422);
   U3043 : OAI21_X1 port map( B1 => n4394, B2 => n4186, A => n83, ZN => n4187);
   U3044 : INV_X1 port map( A => n4187, ZN => n4219);
   U3045 : MUX2_X1 port map( A => n4396, B => n1050, S => n372, Z => n4188);
   U3046 : INV_X1 port map( A => n4188, ZN => n3423);
   U3047 : MUX2_X1 port map( A => n4398, B => n1088, S => n372, Z => n4189);
   U3048 : INV_X1 port map( A => n4189, ZN => n3424);
   U3049 : MUX2_X1 port map( A => n4400, B => n1124, S => n372, Z => n4190);
   U3050 : INV_X1 port map( A => n4190, ZN => n3425);
   U3051 : MUX2_X1 port map( A => n4402, B => n1160, S => n372, Z => n4191);
   U3052 : INV_X1 port map( A => n4191, ZN => n3426);
   U3053 : MUX2_X1 port map( A => n4404, B => n1196, S => n372, Z => n4192);
   U3054 : INV_X1 port map( A => n4192, ZN => n3427);
   U3055 : MUX2_X1 port map( A => n4406, B => n1232, S => n372, Z => n4193);
   U3056 : INV_X1 port map( A => n4193, ZN => n3428);
   U3057 : MUX2_X1 port map( A => n4408, B => n1268, S => n372, Z => n4194);
   U3058 : INV_X1 port map( A => n4194, ZN => n3429);
   U3059 : MUX2_X1 port map( A => n4410, B => n1304, S => n372, Z => n4195);
   U3060 : INV_X1 port map( A => n4195, ZN => n3430);
   U3061 : MUX2_X1 port map( A => n4412, B => n1340, S => n372, Z => n4196);
   U3062 : INV_X1 port map( A => n4196, ZN => n3431);
   U3063 : MUX2_X1 port map( A => n4414, B => n1375, S => n372, Z => n4197);
   U3064 : INV_X1 port map( A => n4197, ZN => n3432);
   U3065 : MUX2_X1 port map( A => n4416, B => n1410, S => n372, Z => n4198);
   U3066 : INV_X1 port map( A => n4198, ZN => n3433);
   U3067 : MUX2_X1 port map( A => n4418, B => n1445, S => n372, Z => n4199);
   U3068 : INV_X1 port map( A => n4199, ZN => n3434);
   U3069 : MUX2_X1 port map( A => n4420, B => n1480, S => n373, Z => n4200);
   U3070 : INV_X1 port map( A => n4200, ZN => n3435);
   U3071 : MUX2_X1 port map( A => n4422, B => n1515, S => n373, Z => n4201);
   U3072 : INV_X1 port map( A => n4201, ZN => n3436);
   U3073 : MUX2_X1 port map( A => n4424, B => n1551, S => n373, Z => n4202);
   U3074 : INV_X1 port map( A => n4202, ZN => n3437);
   U3075 : MUX2_X1 port map( A => n4426, B => n1586, S => n373, Z => n4203);
   U3076 : INV_X1 port map( A => n4203, ZN => n3438);
   U3077 : MUX2_X1 port map( A => n4428, B => n1621, S => n373, Z => n4204);
   U3078 : INV_X1 port map( A => n4204, ZN => n3439);
   U3079 : MUX2_X1 port map( A => n4430, B => n1657, S => n373, Z => n4205);
   U3080 : INV_X1 port map( A => n4205, ZN => n3440);
   U3081 : MUX2_X1 port map( A => n4432, B => n1693, S => n373, Z => n4206);
   U3082 : INV_X1 port map( A => n4206, ZN => n3441);
   U3083 : MUX2_X1 port map( A => n4434, B => n1728, S => n373, Z => n4207);
   U3084 : INV_X1 port map( A => n4207, ZN => n3442);
   U3085 : MUX2_X1 port map( A => n4436, B => n1764, S => n373, Z => n4208);
   U3086 : INV_X1 port map( A => n4208, ZN => n3443);
   U3087 : MUX2_X1 port map( A => n4438, B => n1800, S => n373, Z => n4209);
   U3088 : INV_X1 port map( A => n4209, ZN => n3444);
   U3089 : MUX2_X1 port map( A => n4440, B => n1836, S => n373, Z => n4210);
   U3090 : INV_X1 port map( A => n4210, ZN => n3445);
   U3091 : MUX2_X1 port map( A => n4442, B => n1872, S => n373, Z => n4211);
   U3092 : INV_X1 port map( A => n4211, ZN => n3446);
   U3093 : MUX2_X1 port map( A => n4444, B => n1908, S => n374, Z => n4212);
   U3094 : INV_X1 port map( A => n4212, ZN => n3447);
   U3095 : MUX2_X1 port map( A => n4446, B => n1944, S => n374, Z => n4213);
   U3096 : INV_X1 port map( A => n4213, ZN => n3448);
   U3097 : MUX2_X1 port map( A => n4448, B => n1979, S => n374, Z => n4214);
   U3098 : INV_X1 port map( A => n4214, ZN => n3449);
   U3099 : MUX2_X1 port map( A => n4450, B => n2014, S => n374, Z => n4215);
   U3100 : INV_X1 port map( A => n4215, ZN => n3450);
   U3101 : MUX2_X1 port map( A => n4452, B => n2050, S => n374, Z => n4216);
   U3102 : INV_X1 port map( A => n4216, ZN => n3451);
   U3103 : MUX2_X1 port map( A => n4454, B => n2086, S => n374, Z => n4217);
   U3104 : INV_X1 port map( A => n4217, ZN => n3452);
   U3105 : MUX2_X1 port map( A => n4456, B => n2122, S => n374, Z => n4218);
   U3106 : INV_X1 port map( A => n4218, ZN => n3453);
   U3107 : MUX2_X1 port map( A => n4459, B => n2163, S => n374, Z => n4220);
   U3108 : INV_X1 port map( A => n4220, ZN => n3454);
   U3109 : OAI21_X1 port map( B1 => n4394, B2 => n4221, A => n83, ZN => n4222);
   U3110 : INV_X1 port map( A => n4222, ZN => n4254);
   U3111 : MUX2_X1 port map( A => n4396, B => n1049, S => n375, Z => n4223);
   U3112 : INV_X1 port map( A => n4223, ZN => n3455);
   U3113 : MUX2_X1 port map( A => n4398, B => n1087, S => n375, Z => n4224);
   U3114 : INV_X1 port map( A => n4224, ZN => n3456);
   U3115 : MUX2_X1 port map( A => n4400, B => n1123, S => n375, Z => n4225);
   U3116 : INV_X1 port map( A => n4225, ZN => n3457);
   U3117 : MUX2_X1 port map( A => n4402, B => n1159, S => n375, Z => n4226);
   U3118 : INV_X1 port map( A => n4226, ZN => n3458);
   U3119 : MUX2_X1 port map( A => n4404, B => n1195, S => n375, Z => n4227);
   U3120 : INV_X1 port map( A => n4227, ZN => n3459);
   U3121 : MUX2_X1 port map( A => n4406, B => n1231, S => n375, Z => n4228);
   U3122 : INV_X1 port map( A => n4228, ZN => n3460);
   U3123 : MUX2_X1 port map( A => n4408, B => n1267, S => n375, Z => n4229);
   U3124 : INV_X1 port map( A => n4229, ZN => n3461);
   U3125 : MUX2_X1 port map( A => n4410, B => n1303, S => n375, Z => n4230);
   U3126 : INV_X1 port map( A => n4230, ZN => n3462);
   U3127 : MUX2_X1 port map( A => n4412, B => n1339, S => n375, Z => n4231);
   U3128 : INV_X1 port map( A => n4231, ZN => n3463);
   U3129 : MUX2_X1 port map( A => n4414, B => n1374, S => n375, Z => n4232);
   U3130 : INV_X1 port map( A => n4232, ZN => n3464);
   U3131 : MUX2_X1 port map( A => n4416, B => n1409, S => n375, Z => n4233);
   U3132 : INV_X1 port map( A => n4233, ZN => n3465);
   U3133 : MUX2_X1 port map( A => n4418, B => n1444, S => n375, Z => n4234);
   U3134 : INV_X1 port map( A => n4234, ZN => n3466);
   U3135 : MUX2_X1 port map( A => n4420, B => n1479, S => n376, Z => n4235);
   U3136 : INV_X1 port map( A => n4235, ZN => n3467);
   U3137 : MUX2_X1 port map( A => n4422, B => n1514, S => n376, Z => n4236);
   U3138 : INV_X1 port map( A => n4236, ZN => n3468);
   U3139 : MUX2_X1 port map( A => n4424, B => n1550, S => n376, Z => n4237);
   U3140 : INV_X1 port map( A => n4237, ZN => n3469);
   U3141 : MUX2_X1 port map( A => n4426, B => n1585, S => n376, Z => n4238);
   U3142 : INV_X1 port map( A => n4238, ZN => n3470);
   U3143 : MUX2_X1 port map( A => n4428, B => n1620, S => n376, Z => n4239);
   U3144 : INV_X1 port map( A => n4239, ZN => n3471);
   U3145 : MUX2_X1 port map( A => n4430, B => n1656, S => n376, Z => n4240);
   U3146 : INV_X1 port map( A => n4240, ZN => n3472);
   U3147 : MUX2_X1 port map( A => n4432, B => n1692, S => n376, Z => n4241);
   U3148 : INV_X1 port map( A => n4241, ZN => n3473);
   U3149 : MUX2_X1 port map( A => n4434, B => n1727, S => n376, Z => n4242);
   U3150 : INV_X1 port map( A => n4242, ZN => n3474);
   U3151 : MUX2_X1 port map( A => n4436, B => n1763, S => n376, Z => n4243);
   U3152 : INV_X1 port map( A => n4243, ZN => n3475);
   U3153 : MUX2_X1 port map( A => n4438, B => n1799, S => n376, Z => n4244);
   U3154 : INV_X1 port map( A => n4244, ZN => n3476);
   U3155 : MUX2_X1 port map( A => n4440, B => n1835, S => n376, Z => n4245);
   U3156 : INV_X1 port map( A => n4245, ZN => n3477);
   U3157 : MUX2_X1 port map( A => n4442, B => n1871, S => n376, Z => n4246);
   U3158 : INV_X1 port map( A => n4246, ZN => n3478);
   U3159 : MUX2_X1 port map( A => n4444, B => n1907, S => n377, Z => n4247);
   U3160 : INV_X1 port map( A => n4247, ZN => n3479);
   U3161 : MUX2_X1 port map( A => n4446, B => n1943, S => n377, Z => n4248);
   U3162 : INV_X1 port map( A => n4248, ZN => n3480);
   U3163 : MUX2_X1 port map( A => n4448, B => n1978, S => n377, Z => n4249);
   U3164 : INV_X1 port map( A => n4249, ZN => n3481);
   U3165 : MUX2_X1 port map( A => n4450, B => n2013, S => n377, Z => n4250);
   U3166 : INV_X1 port map( A => n4250, ZN => n3482);
   U3167 : MUX2_X1 port map( A => n4452, B => n2049, S => n377, Z => n4251);
   U3168 : INV_X1 port map( A => n4251, ZN => n3483);
   U3169 : MUX2_X1 port map( A => n4454, B => n2085, S => n377, Z => n4252);
   U3170 : INV_X1 port map( A => n4252, ZN => n3484);
   U3171 : MUX2_X1 port map( A => n4456, B => n2121, S => n377, Z => n4253);
   U3172 : INV_X1 port map( A => n4253, ZN => n3485);
   U3173 : MUX2_X1 port map( A => n4459, B => n2161, S => n377, Z => n4255);
   U3174 : INV_X1 port map( A => n4255, ZN => n3486);
   U3175 : OAI21_X1 port map( B1 => n4394, B2 => n4256, A => n83, ZN => n4257);
   U3176 : INV_X1 port map( A => n4257, ZN => n4289);
   U3177 : MUX2_X1 port map( A => n4294, B => n4258, S => n378, Z => n3487);
   U3178 : MUX2_X1 port map( A => n4296, B => n4259, S => n378, Z => n3488);
   U3179 : MUX2_X1 port map( A => n4298, B => n4260, S => n378, Z => n3489);
   U3180 : MUX2_X1 port map( A => n4300, B => n4261, S => n378, Z => n3490);
   U3181 : MUX2_X1 port map( A => n4302, B => n4262, S => n378, Z => n3491);
   U3182 : MUX2_X1 port map( A => n4304, B => n4263, S => n378, Z => n3492);
   U3183 : MUX2_X1 port map( A => n4306, B => n4264, S => n378, Z => n3493);
   U3184 : MUX2_X1 port map( A => n4308, B => n4265, S => n378, Z => n3494);
   U3185 : MUX2_X1 port map( A => n4310, B => n4266, S => n378, Z => n3495);
   U3186 : MUX2_X1 port map( A => n4312, B => n4267, S => n378, Z => n3496);
   U3187 : MUX2_X1 port map( A => n4314, B => n4268, S => n378, Z => n3497);
   U3188 : MUX2_X1 port map( A => n4316, B => n4269, S => n378, Z => n3498);
   U3189 : MUX2_X1 port map( A => n4318, B => n4270, S => n379, Z => n3499);
   U3190 : MUX2_X1 port map( A => n4320, B => n4271, S => n379, Z => n3500);
   U3191 : MUX2_X1 port map( A => n4322, B => n4272, S => n379, Z => n3501);
   U3192 : MUX2_X1 port map( A => n4324, B => n4273, S => n379, Z => n3502);
   U3193 : MUX2_X1 port map( A => n4326, B => n4274, S => n379, Z => n3503);
   U3194 : MUX2_X1 port map( A => n4328, B => n4275, S => n379, Z => n3504);
   U3195 : MUX2_X1 port map( A => n4330, B => n4276, S => n379, Z => n3505);
   U3196 : MUX2_X1 port map( A => n4332, B => n4277, S => n379, Z => n3506);
   U3197 : MUX2_X1 port map( A => n4334, B => n4278, S => n379, Z => n3507);
   U3198 : MUX2_X1 port map( A => n4336, B => n4279, S => n379, Z => n3508);
   U3199 : MUX2_X1 port map( A => n4338, B => n4280, S => n379, Z => n3509);
   U3200 : MUX2_X1 port map( A => n4340, B => n4281, S => n379, Z => n3510);
   U3201 : MUX2_X1 port map( A => n4342, B => n4282, S => n380, Z => n3511);
   U3202 : MUX2_X1 port map( A => n4344, B => n4283, S => n380, Z => n3512);
   U3203 : MUX2_X1 port map( A => n4346, B => n4284, S => n380, Z => n3513);
   U3204 : MUX2_X1 port map( A => n4348, B => n4285, S => n380, Z => n3514);
   U3205 : MUX2_X1 port map( A => n4350, B => n4286, S => n380, Z => n3515);
   U3206 : MUX2_X1 port map( A => n4352, B => n4287, S => n380, Z => n3516);
   U3207 : MUX2_X1 port map( A => n4354, B => n4288, S => n380, Z => n3517);
   U3208 : MUX2_X1 port map( A => n4357, B => n4290, S => n380, Z => n3518);
   U3209 : OAI21_X1 port map( B1 => n4394, B2 => n4291, A => n83, ZN => n4292);
   U3210 : INV_X1 port map( A => n4292, ZN => n4355);
   U3211 : MUX2_X1 port map( A => n4294, B => n4293, S => n381, Z => n3519);
   U3212 : MUX2_X1 port map( A => n4296, B => n4295, S => n381, Z => n3520);
   U3213 : MUX2_X1 port map( A => n4298, B => n4297, S => n381, Z => n3521);
   U3214 : MUX2_X1 port map( A => n4300, B => n4299, S => n381, Z => n3522);
   U3215 : MUX2_X1 port map( A => n4302, B => n4301, S => n381, Z => n3523);
   U3216 : MUX2_X1 port map( A => n4304, B => n4303, S => n381, Z => n3524);
   U3217 : MUX2_X1 port map( A => n4306, B => n4305, S => n381, Z => n3525);
   U3218 : MUX2_X1 port map( A => n4308, B => n4307, S => n381, Z => n3526);
   U3219 : MUX2_X1 port map( A => n4310, B => n4309, S => n381, Z => n3527);
   U3220 : MUX2_X1 port map( A => n4312, B => n4311, S => n381, Z => n3528);
   U3221 : MUX2_X1 port map( A => n4314, B => n4313, S => n381, Z => n3529);
   U3222 : MUX2_X1 port map( A => n4316, B => n4315, S => n381, Z => n3530);
   U3223 : MUX2_X1 port map( A => n4318, B => n4317, S => n382, Z => n3531);
   U3224 : MUX2_X1 port map( A => n4320, B => n4319, S => n382, Z => n3532);
   U3225 : MUX2_X1 port map( A => n4322, B => n4321, S => n382, Z => n3533);
   U3226 : MUX2_X1 port map( A => n4324, B => n4323, S => n382, Z => n3534);
   U3227 : MUX2_X1 port map( A => n4326, B => n4325, S => n382, Z => n3535);
   U3228 : MUX2_X1 port map( A => n4328, B => n4327, S => n382, Z => n3536);
   U3229 : MUX2_X1 port map( A => n4330, B => n4329, S => n382, Z => n3537);
   U3230 : MUX2_X1 port map( A => n4332, B => n4331, S => n382, Z => n3538);
   U3231 : MUX2_X1 port map( A => n4334, B => n4333, S => n382, Z => n3539);
   U3232 : MUX2_X1 port map( A => n4336, B => n4335, S => n382, Z => n3540);
   U3233 : MUX2_X1 port map( A => n4338, B => n4337, S => n382, Z => n3541);
   U3234 : MUX2_X1 port map( A => n4340, B => n4339, S => n382, Z => n3542);
   U3235 : MUX2_X1 port map( A => n4342, B => n4341, S => n383, Z => n3543);
   U3236 : MUX2_X1 port map( A => n4344, B => n4343, S => n383, Z => n3544);
   U3237 : MUX2_X1 port map( A => n4346, B => n4345, S => n383, Z => n3545);
   U3238 : MUX2_X1 port map( A => n4348, B => n4347, S => n383, Z => n3546);
   U3239 : MUX2_X1 port map( A => n4350, B => n4349, S => n383, Z => n3547);
   U3240 : MUX2_X1 port map( A => n4352, B => n4351, S => n383, Z => n3548);
   U3241 : MUX2_X1 port map( A => n4354, B => n4353, S => n383, Z => n3549);
   U3242 : MUX2_X1 port map( A => n4357, B => n4356, S => n383, Z => n3550);
   U3243 : OAI21_X1 port map( B1 => n4394, B2 => n4358, A => n83, ZN => n4359);
   U3244 : INV_X1 port map( A => n4359, ZN => n4391);
   U3245 : MUX2_X1 port map( A => n4396, B => n1053, S => n384, Z => n4360);
   U3246 : INV_X1 port map( A => n4360, ZN => n3551);
   U3247 : MUX2_X1 port map( A => n4398, B => n1091, S => n384, Z => n4361);
   U3248 : INV_X1 port map( A => n4361, ZN => n3552);
   U3249 : MUX2_X1 port map( A => n4400, B => n1127, S => n384, Z => n4362);
   U3250 : INV_X1 port map( A => n4362, ZN => n3553);
   U3251 : MUX2_X1 port map( A => n4402, B => n1163, S => n384, Z => n4363);
   U3252 : INV_X1 port map( A => n4363, ZN => n3554);
   U3253 : MUX2_X1 port map( A => n4404, B => n1199, S => n384, Z => n4364);
   U3254 : INV_X1 port map( A => n4364, ZN => n3555);
   U3255 : MUX2_X1 port map( A => n4406, B => n1235, S => n384, Z => n4365);
   U3256 : INV_X1 port map( A => n4365, ZN => n3556);
   U3257 : MUX2_X1 port map( A => n4408, B => n1271, S => n384, Z => n4366);
   U3258 : INV_X1 port map( A => n4366, ZN => n3557);
   U3259 : MUX2_X1 port map( A => n4410, B => n1307, S => n384, Z => n4367);
   U3260 : INV_X1 port map( A => n4367, ZN => n3558);
   U3261 : MUX2_X1 port map( A => n4412, B => n1343, S => n384, Z => n4368);
   U3262 : INV_X1 port map( A => n4368, ZN => n3559);
   U3263 : MUX2_X1 port map( A => n4414, B => n1378, S => n384, Z => n4369);
   U3264 : INV_X1 port map( A => n4369, ZN => n3560);
   U3265 : MUX2_X1 port map( A => n4416, B => n1413, S => n384, Z => n4370);
   U3266 : INV_X1 port map( A => n4370, ZN => n3561);
   U3267 : MUX2_X1 port map( A => n4418, B => n1448, S => n384, Z => n4371);
   U3268 : INV_X1 port map( A => n4371, ZN => n3562);
   U3269 : MUX2_X1 port map( A => n4420, B => n1483, S => n385, Z => n4372);
   U3270 : INV_X1 port map( A => n4372, ZN => n3563);
   U3271 : MUX2_X1 port map( A => n4422, B => n1518, S => n385, Z => n4373);
   U3272 : INV_X1 port map( A => n4373, ZN => n3564);
   U3273 : MUX2_X1 port map( A => n4424, B => n1554, S => n385, Z => n4374);
   U3274 : INV_X1 port map( A => n4374, ZN => n3565);
   U3275 : MUX2_X1 port map( A => n4426, B => n1589, S => n385, Z => n4375);
   U3276 : INV_X1 port map( A => n4375, ZN => n3566);
   U3277 : MUX2_X1 port map( A => n4428, B => n1624, S => n385, Z => n4376);
   U3278 : INV_X1 port map( A => n4376, ZN => n3567);
   U3279 : MUX2_X1 port map( A => n4430, B => n1660, S => n385, Z => n4377);
   U3280 : INV_X1 port map( A => n4377, ZN => n3568);
   U3281 : MUX2_X1 port map( A => n4432, B => n1696, S => n385, Z => n4378);
   U3282 : INV_X1 port map( A => n4378, ZN => n3569);
   U3283 : MUX2_X1 port map( A => n4434, B => n1731, S => n385, Z => n4379);
   U3284 : INV_X1 port map( A => n4379, ZN => n3570);
   U3285 : MUX2_X1 port map( A => n4436, B => n1767, S => n385, Z => n4380);
   U3286 : INV_X1 port map( A => n4380, ZN => n3571);
   U3287 : MUX2_X1 port map( A => n4438, B => n1803, S => n385, Z => n4381);
   U3288 : INV_X1 port map( A => n4381, ZN => n3572);
   U3289 : MUX2_X1 port map( A => n4440, B => n1839, S => n385, Z => n4382);
   U3290 : INV_X1 port map( A => n4382, ZN => n3573);
   U3291 : MUX2_X1 port map( A => n4442, B => n1875, S => n385, Z => n4383);
   U3292 : INV_X1 port map( A => n4383, ZN => n3574);
   U3293 : MUX2_X1 port map( A => n4444, B => n1911, S => n386, Z => n4384);
   U3294 : INV_X1 port map( A => n4384, ZN => n3575);
   U3295 : MUX2_X1 port map( A => n4446, B => n1947, S => n386, Z => n4385);
   U3296 : INV_X1 port map( A => n4385, ZN => n3576);
   U3297 : MUX2_X1 port map( A => n4448, B => n1982, S => n386, Z => n4386);
   U3298 : INV_X1 port map( A => n4386, ZN => n3577);
   U3299 : MUX2_X1 port map( A => n4450, B => n2017, S => n386, Z => n4387);
   U3300 : INV_X1 port map( A => n4387, ZN => n3578);
   U3301 : MUX2_X1 port map( A => n4452, B => n2053, S => n386, Z => n4388);
   U3302 : INV_X1 port map( A => n4388, ZN => n3579);
   U3303 : MUX2_X1 port map( A => n4454, B => n2089, S => n386, Z => n4389);
   U3304 : INV_X1 port map( A => n4389, ZN => n3580);
   U3305 : MUX2_X1 port map( A => n4456, B => n2125, S => n386, Z => n4390);
   U3306 : INV_X1 port map( A => n4390, ZN => n3581);
   U3307 : MUX2_X1 port map( A => n4459, B => n2168, S => n386, Z => n4392);
   U3308 : INV_X1 port map( A => n4392, ZN => n3582);
   U3309 : OAI21_X1 port map( B1 => n4394, B2 => n4393, A => n84, ZN => n4395);
   U3310 : INV_X1 port map( A => n4395, ZN => n4458);
   U3311 : MUX2_X1 port map( A => n4396, B => n1052, S => n387, Z => n4397);
   U3312 : INV_X1 port map( A => n4397, ZN => n3583);
   U3313 : MUX2_X1 port map( A => n4398, B => n1090, S => n387, Z => n4399);
   U3314 : INV_X1 port map( A => n4399, ZN => n3584);
   U3315 : MUX2_X1 port map( A => n4400, B => n1126, S => n387, Z => n4401);
   U3316 : INV_X1 port map( A => n4401, ZN => n3585);
   U3317 : MUX2_X1 port map( A => n4402, B => n1162, S => n387, Z => n4403);
   U3318 : INV_X1 port map( A => n4403, ZN => n3586);
   U3319 : MUX2_X1 port map( A => n4404, B => n1198, S => n387, Z => n4405);
   U3320 : INV_X1 port map( A => n4405, ZN => n3587);
   U3321 : MUX2_X1 port map( A => n4406, B => n1234, S => n387, Z => n4407);
   U3322 : INV_X1 port map( A => n4407, ZN => n3588);
   U3323 : MUX2_X1 port map( A => n4408, B => n1270, S => n387, Z => n4409);
   U3324 : INV_X1 port map( A => n4409, ZN => n3589);
   U3325 : MUX2_X1 port map( A => n4410, B => n1306, S => n387, Z => n4411);
   U3326 : INV_X1 port map( A => n4411, ZN => n3590);
   U3327 : MUX2_X1 port map( A => n4412, B => n1342, S => n387, Z => n4413);
   U3328 : INV_X1 port map( A => n4413, ZN => n3591);
   U3329 : MUX2_X1 port map( A => n4414, B => n1377, S => n387, Z => n4415);
   U3330 : INV_X1 port map( A => n4415, ZN => n3592);
   U3331 : MUX2_X1 port map( A => n4416, B => n1412, S => n387, Z => n4417);
   U3332 : INV_X1 port map( A => n4417, ZN => n3593);
   U3333 : MUX2_X1 port map( A => n4418, B => n1447, S => n387, Z => n4419);
   U3334 : INV_X1 port map( A => n4419, ZN => n3594);
   U3335 : MUX2_X1 port map( A => n4420, B => n1482, S => n388, Z => n4421);
   U3336 : INV_X1 port map( A => n4421, ZN => n3595);
   U3337 : MUX2_X1 port map( A => n4422, B => n1517, S => n388, Z => n4423);
   U3338 : INV_X1 port map( A => n4423, ZN => n3596);
   U3339 : MUX2_X1 port map( A => n4424, B => n1553, S => n388, Z => n4425);
   U3340 : INV_X1 port map( A => n4425, ZN => n3597);
   U3341 : MUX2_X1 port map( A => n4426, B => n1588, S => n388, Z => n4427);
   U3342 : INV_X1 port map( A => n4427, ZN => n3598);
   U3343 : MUX2_X1 port map( A => n4428, B => n1623, S => n388, Z => n4429);
   U3344 : INV_X1 port map( A => n4429, ZN => n3599);
   U3345 : MUX2_X1 port map( A => n4430, B => n1659, S => n388, Z => n4431);
   U3346 : INV_X1 port map( A => n4431, ZN => n3600);
   U3347 : MUX2_X1 port map( A => n4432, B => n1695, S => n388, Z => n4433);
   U3348 : INV_X1 port map( A => n4433, ZN => n3601);
   U3349 : MUX2_X1 port map( A => n4434, B => n1730, S => n388, Z => n4435);
   U3350 : INV_X1 port map( A => n4435, ZN => n3602);
   U3351 : MUX2_X1 port map( A => n4436, B => n1766, S => n388, Z => n4437);
   U3352 : INV_X1 port map( A => n4437, ZN => n3603);
   U3353 : MUX2_X1 port map( A => n4438, B => n1802, S => n388, Z => n4439);
   U3354 : INV_X1 port map( A => n4439, ZN => n3604);
   U3355 : MUX2_X1 port map( A => n4440, B => n1838, S => n388, Z => n4441);
   U3356 : INV_X1 port map( A => n4441, ZN => n3605);
   U3357 : MUX2_X1 port map( A => n4442, B => n1874, S => n388, Z => n4443);
   U3358 : INV_X1 port map( A => n4443, ZN => n3606);
   U3359 : MUX2_X1 port map( A => n4444, B => n1910, S => n389, Z => n4445);
   U3360 : INV_X1 port map( A => n4445, ZN => n3607);
   U3361 : MUX2_X1 port map( A => n4446, B => n1946, S => n389, Z => n4447);
   U3362 : INV_X1 port map( A => n4447, ZN => n3608);
   U3363 : MUX2_X1 port map( A => n4448, B => n1981, S => n389, Z => n4449);
   U3364 : INV_X1 port map( A => n4449, ZN => n3609);
   U3365 : MUX2_X1 port map( A => n4450, B => n2016, S => n389, Z => n4451);
   U3366 : INV_X1 port map( A => n4451, ZN => n3610);
   U3367 : MUX2_X1 port map( A => n4452, B => n2052, S => n389, Z => n4453);
   U3368 : INV_X1 port map( A => n4453, ZN => n3611);
   U3369 : MUX2_X1 port map( A => n4454, B => n2088, S => n389, Z => n4455);
   U3370 : INV_X1 port map( A => n4455, ZN => n3612);
   U3371 : MUX2_X1 port map( A => n4456, B => n2124, S => n389, Z => n4457);
   U3372 : INV_X1 port map( A => n4457, ZN => n3613);
   U3373 : MUX2_X1 port map( A => n4459, B => n2166, S => n389, Z => n4460);
   U3374 : INV_X1 port map( A => n4460, ZN => n3614);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => OUT2(10), QN
                           => n20);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => OUT2(9), QN 
                           => n590);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => OUT2(8), QN 
                           => n570);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => OUT2(7), QN 
                           => n8);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => OUT2(6), QN 
                           => n7);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => OUT2(5), QN 
                           => n512);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => OUT2(4), QN 
                           => n492);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => OUT2(3), QN 
                           => n472);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => OUT2(2), QN 
                           => n88);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => OUT2(1), QN 
                           => n89);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2527, CK => CLK, Q => OUT2(0), QN 
                           => n414);
   OUT1_reg_31_inst : DFF_X1 port map( D => n2590, CK => CLK, Q => OUT1(31), QN
                           => n2202);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2589, CK => CLK, Q => OUT1(30), QN
                           => n2150);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2588, CK => CLK, Q => OUT1(29), QN
                           => n2114);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2587, CK => CLK, Q => OUT1(28), QN
                           => n2078);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2586, CK => CLK, Q => OUT1(27), QN
                           => n2042);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2585, CK => CLK, Q => OUT1(26), QN
                           => n5);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2584, CK => CLK, Q => OUT1(25), QN
                           => n6);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2583, CK => CLK, Q => OUT1(24), QN
                           => n1936);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => OUT2(11), QN
                           => n9);
   OUT2_reg_31_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => OUT2(31), QN
                           => n1038);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => OUT2(30), QN
                           => n1002);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => OUT2(29), QN
                           => n982);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => OUT2(28), QN
                           => n962);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => OUT2(27), QN
                           => n942);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => OUT2(26), QN
                           => n12);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => OUT2(25), QN
                           => n903);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => OUT2(24), QN
                           => n14);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => OUT1(10), QN
                           => n26);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => OUT1(9), QN 
                           => n23);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => OUT1(8), QN 
                           => n19);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => OUT1(7), QN 
                           => n1332);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => OUT1(6), QN 
                           => n1296);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_N32 is

   port( CURR_ADDR : in std_logic_vector (31 downto 0);  NEXT_ADDR : out 
         std_logic_vector (31 downto 0));

end ADDER_N32;

architecture SYN_BEHAVIOR of ADDER_N32 is

   component ADDER_N32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n3, n_2185 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '1';
   n3 <= '0';
   add_26 : ADDER_N32_DW01_add_0 port map( A(31) => CURR_ADDR(31), A(30) => 
                           CURR_ADDR(30), A(29) => CURR_ADDR(29), A(28) => 
                           CURR_ADDR(28), A(27) => CURR_ADDR(27), A(26) => 
                           CURR_ADDR(26), A(25) => CURR_ADDR(25), A(24) => 
                           CURR_ADDR(24), A(23) => CURR_ADDR(23), A(22) => 
                           CURR_ADDR(22), A(21) => CURR_ADDR(21), A(20) => 
                           CURR_ADDR(20), A(19) => CURR_ADDR(19), A(18) => 
                           CURR_ADDR(18), A(17) => CURR_ADDR(17), A(16) => 
                           CURR_ADDR(16), A(15) => CURR_ADDR(15), A(14) => 
                           CURR_ADDR(14), A(13) => CURR_ADDR(13), A(12) => 
                           CURR_ADDR(12), A(11) => CURR_ADDR(11), A(10) => 
                           CURR_ADDR(10), A(9) => CURR_ADDR(9), A(8) => 
                           CURR_ADDR(8), A(7) => CURR_ADDR(7), A(6) => 
                           CURR_ADDR(6), A(5) => CURR_ADDR(5), A(4) => 
                           CURR_ADDR(4), A(3) => CURR_ADDR(3), A(2) => 
                           CURR_ADDR(2), A(1) => CURR_ADDR(1), A(0) => 
                           CURR_ADDR(0), B(31) => n1, B(30) => n1, B(29) => n1,
                           B(28) => n1, B(27) => n1, B(26) => n1, B(25) => n1, 
                           B(24) => n1, B(23) => n1, B(22) => n1, B(21) => n1, 
                           B(20) => n1, B(19) => n1, B(18) => n1, B(17) => n1, 
                           B(16) => n1, B(15) => n1, B(14) => n1, B(13) => n1, 
                           B(12) => n1, B(11) => n1, B(10) => n1, B(9) => n1, 
                           B(8) => n1, B(7) => n1, B(6) => n1, B(5) => n1, B(4)
                           => n1, B(3) => n1, B(2) => n2, B(1) => n1, B(0) => 
                           n1, CI => n3, SUM(31) => NEXT_ADDR(31), SUM(30) => 
                           NEXT_ADDR(30), SUM(29) => NEXT_ADDR(29), SUM(28) => 
                           NEXT_ADDR(28), SUM(27) => NEXT_ADDR(27), SUM(26) => 
                           NEXT_ADDR(26), SUM(25) => NEXT_ADDR(25), SUM(24) => 
                           NEXT_ADDR(24), SUM(23) => NEXT_ADDR(23), SUM(22) => 
                           NEXT_ADDR(22), SUM(21) => NEXT_ADDR(21), SUM(20) => 
                           NEXT_ADDR(20), SUM(19) => NEXT_ADDR(19), SUM(18) => 
                           NEXT_ADDR(18), SUM(17) => NEXT_ADDR(17), SUM(16) => 
                           NEXT_ADDR(16), SUM(15) => NEXT_ADDR(15), SUM(14) => 
                           NEXT_ADDR(14), SUM(13) => NEXT_ADDR(13), SUM(12) => 
                           NEXT_ADDR(12), SUM(11) => NEXT_ADDR(11), SUM(10) => 
                           NEXT_ADDR(10), SUM(9) => NEXT_ADDR(9), SUM(8) => 
                           NEXT_ADDR(8), SUM(7) => NEXT_ADDR(7), SUM(6) => 
                           NEXT_ADDR(6), SUM(5) => NEXT_ADDR(5), SUM(4) => 
                           NEXT_ADDR(4), SUM(3) => NEXT_ADDR(3), SUM(2) => 
                           NEXT_ADDR(2), SUM(1) => NEXT_ADDR(1), SUM(0) => 
                           NEXT_ADDR(0), CO => n_2185);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT5_1 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_GENERIC_NBIT5_1;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n12, n13, n14, n15, n16 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n12, ZN => Y(0));
   U2 : AOI22_X1 port map( A1 => A(0), A2 => n6, B1 => B(0), B2 => SEL, ZN => 
                           n12);
   U3 : INV_X1 port map( A => n13, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n6, B1 => B(1), B2 => SEL, ZN => 
                           n13);
   U5 : INV_X1 port map( A => n14, ZN => Y(2));
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n6, B1 => B(2), B2 => SEL, ZN => 
                           n14);
   U7 : INV_X1 port map( A => n15, ZN => Y(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n6, B1 => B(3), B2 => SEL, ZN => 
                           n15);
   U9 : INV_X1 port map( A => n16, ZN => Y(4));
   U10 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => SEL, B2 => B(4), ZN => 
                           n16);
   U11 : INV_X1 port map( A => SEL, ZN => n6);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_2;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_3;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal net50426, n1 : std_logic;

begin
   
   U1 : MUX2_X2 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U2 : MUX2_X2 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U3 : MUX2_X2 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U4 : MUX2_X2 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U5 : MUX2_X2 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U6 : MUX2_X2 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U7 : MUX2_X2 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U8 : MUX2_X2 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X2 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U10 : MUX2_X2 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U11 : MUX2_X2 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U12 : MUX2_X2 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U13 : MUX2_X2 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U14 : MUX2_X2 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : INV_X1 port map( A => n1, ZN => Y(2));
   U16 : MUX2_X2 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U17 : MUX2_X2 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U18 : MUX2_X2 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U19 : MUX2_X2 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U20 : MUX2_X2 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U21 : MUX2_X2 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U22 : MUX2_X2 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U23 : MUX2_X2 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U24 : MUX2_X2 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U25 : MUX2_X2 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U26 : INV_X1 port map( A => SEL, ZN => net50426);
   U27 : AOI22_X1 port map( A1 => A(2), A2 => net50426, B1 => B(2), B2 => SEL, 
                           ZN => n1);
   U28 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U29 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U30 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U31 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U32 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U33 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U34 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_4;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Y(1));
   U2 : MUX2_X2 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U3 : INV_X2 port map( A => n1, ZN => Y(0));
   U4 : MUX2_X2 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U5 : MUX2_X2 port map( A => B(5), B => A(5), S => n4, Z => Y(5));
   U6 : MUX2_X2 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U7 : MUX2_X2 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U8 : MUX2_X2 port map( A => B(12), B => A(12), S => n4, Z => Y(12));
   U9 : INV_X1 port map( A => n3, ZN => Y(2));
   U10 : MUX2_X2 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U11 : MUX2_X2 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U12 : MUX2_X2 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U13 : MUX2_X2 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U14 : INV_X1 port map( A => n5, ZN => Y(8));
   U15 : MUX2_X2 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U16 : MUX2_X2 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U17 : MUX2_X2 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U18 : MUX2_X2 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U19 : MUX2_X2 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U20 : MUX2_X2 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U21 : MUX2_X2 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U22 : MUX2_X2 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U23 : MUX2_X2 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U24 : MUX2_X2 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U25 : MUX2_X2 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U26 : MUX2_X2 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U27 : MUX2_X2 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U28 : MUX2_X2 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U29 : MUX2_X2 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U30 : MUX2_X2 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U31 : MUX2_X2 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U32 : INV_X1 port map( A => SEL, ZN => n4);
   U33 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => SEL, ZN => 
                           n1);
   U34 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => SEL, ZN => 
                           n2);
   U35 : AOI22_X1 port map( A1 => A(2), A2 => n4, B1 => B(2), B2 => SEL, ZN => 
                           n3);
   U36 : AOI22_X1 port map( A1 => A(8), A2 => n4, B1 => B(8), B2 => SEL, ZN => 
                           n5);
   U37 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT5_0 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_GENERIC_NBIT5_0;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT5_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21 is

   port( A, B, SEL : in std_logic;  Y : out std_logic);

end MUX21;

architecture SYN_BEHAVIOR of MUX21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => SEL, B2 => B, ZN => n3);
   U3 : INV_X1 port map( A => SEL, ZN => n2);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_0;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : BUF_X1 port map( A => SEL, Z => n3);
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U5 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U6 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U7 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U8 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U9 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U11 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U12 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U13 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U14 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U15 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U16 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U17 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U20 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U21 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U22 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U23 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U24 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U26 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U27 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U28 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U29 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U30 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U31 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Y(27));
   U32 : MUX2_X1 port map( A => A(28), B => B(28), S => n3, Z => Y(28));
   U33 : MUX2_X1 port map( A => A(29), B => B(29), S => n3, Z => Y(29));
   U34 : MUX2_X1 port map( A => A(30), B => B(30), S => n3, Z => Y(30));
   U35 : MUX2_X1 port map( A => A(31), B => B(31), S => n3, Z => Y(31));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BRANCHING_UNIT_N32 is

   port( CLK, RST : in std_logic;  Reg_A : in std_logic_vector (31 downto 0);  
         EQ_cond, IS_JUMP : in std_logic;  branch_taken : out std_logic);

end BRANCHING_UNIT_N32;

architecture SYN_BEHAVIOR of BRANCHING_UNIT_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n_2186 :
      std_logic;

begin
   
   branch_taken_reg : DFF_X1 port map( D => n14, CK => CLK, Q => branch_taken, 
                           QN => n_2186);
   U3 : NOR4_X1 port map( A1 => Reg_A(19), A2 => Reg_A(18), A3 => Reg_A(17), A4
                           => Reg_A(16), ZN => n4);
   U4 : NOR4_X1 port map( A1 => Reg_A(23), A2 => Reg_A(22), A3 => Reg_A(21), A4
                           => Reg_A(20), ZN => n3);
   U5 : NOR4_X1 port map( A1 => Reg_A(27), A2 => Reg_A(26), A3 => Reg_A(25), A4
                           => Reg_A(24), ZN => n2);
   U6 : NOR4_X1 port map( A1 => Reg_A(31), A2 => Reg_A(30), A3 => Reg_A(29), A4
                           => Reg_A(28), ZN => n1);
   U7 : NAND4_X1 port map( A1 => n4, A2 => n3, A3 => n2, A4 => n1, ZN => n10);
   U8 : NOR4_X1 port map( A1 => Reg_A(3), A2 => Reg_A(2), A3 => Reg_A(1), A4 =>
                           Reg_A(0), ZN => n8);
   U9 : NOR4_X1 port map( A1 => Reg_A(7), A2 => Reg_A(6), A3 => Reg_A(5), A4 =>
                           Reg_A(4), ZN => n7);
   U10 : NOR4_X1 port map( A1 => Reg_A(11), A2 => Reg_A(10), A3 => Reg_A(9), A4
                           => Reg_A(8), ZN => n6);
   U11 : NOR4_X1 port map( A1 => Reg_A(15), A2 => Reg_A(14), A3 => Reg_A(13), 
                           A4 => Reg_A(12), ZN => n5);
   U12 : NAND4_X1 port map( A1 => n8, A2 => n7, A3 => n6, A4 => n5, ZN => n9);
   U13 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n11);
   U14 : XNOR2_X1 port map( A => EQ_cond, B => n11, ZN => n12);
   U15 : OAI21_X1 port map( B1 => IS_JUMP, B2 => n12, A => RST, ZN => n13);
   U16 : INV_X1 port map( A => n13, ZN => n14);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_1 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_1;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n36, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193,
      n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, 
      n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, 
      n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218 : std_logic;

begin
   DATA_OUT <= ( DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port );
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n9, CK => CLK, Q => 
                           DATA_OUT_31_port, QN => n_2187);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n10, CK => CLK, Q => 
                           DATA_OUT_30_port, QN => n_2188);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n11, CK => CLK, Q => 
                           DATA_OUT_29_port, QN => n_2189);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n12, CK => CLK, Q => 
                           DATA_OUT_28_port, QN => n_2190);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n13, CK => CLK, Q => 
                           DATA_OUT_27_port, QN => n_2191);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n14, CK => CLK, Q => 
                           DATA_OUT_26_port, QN => n_2192);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n15, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_2193);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n16, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n_2194);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n17, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_2195);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n18, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n_2196);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n19, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n_2197);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n20, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_2198);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n21, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_2199);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n22, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_2200);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n23, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_2201);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n24, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n_2202);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n25, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n_2203);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n26, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n_2204);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n27, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n_2205);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n28, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n_2206);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n29, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n_2207);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n30, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n_2208);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n31, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n_2209);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n32, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n_2210);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n33, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n_2211);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n36, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n_2212);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT_5_port, QN => n_2213);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_2214);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_2215);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_2216);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_2217);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_2218);
   U22 : AOI22_X1 port map( A1 => DATA_IN(19), A2 => n7, B1 => DATA_OUT_19_port
                           , B2 => n4, ZN => n86);
   U3 : AOI22_X1 port map( A1 => DATA_IN(0), A2 => n8, B1 => DATA_OUT_0_port, 
                           B2 => n3, ZN => n106);
   U31 : AOI22_X1 port map( A1 => DATA_IN(28), A2 => n6, B1 => DATA_OUT_28_port
                           , B2 => n5, ZN => n77);
   U8 : AOI22_X1 port map( A1 => DATA_IN(5), A2 => n8, B1 => DATA_OUT_5_port, 
                           B2 => n3, ZN => n100);
   U7 : AOI22_X1 port map( A1 => DATA_IN(4), A2 => n8, B1 => DATA_OUT_4_port, 
                           B2 => n3, ZN => n101);
   U6 : AOI22_X1 port map( A1 => DATA_IN(3), A2 => n8, B1 => DATA_OUT_3_port, 
                           B2 => n3, ZN => n102);
   U5 : AOI22_X1 port map( A1 => DATA_IN(2), A2 => n8, B1 => DATA_OUT_2_port, 
                           B2 => n3, ZN => n103);
   U4 : AOI22_X1 port map( A1 => DATA_IN(1), A2 => n8, B1 => DATA_OUT_1_port, 
                           B2 => n3, ZN => n104);
   U10 : AOI22_X1 port map( A1 => DATA_IN(7), A2 => n8, B1 => DATA_OUT_7_port, 
                           B2 => n3, ZN => n98);
   U9 : AOI22_X1 port map( A1 => DATA_IN(6), A2 => n8, B1 => DATA_OUT_6_port, 
                           B2 => n3, ZN => n99);
   U34 : AOI22_X1 port map( A1 => DATA_IN(31), A2 => n6, B1 => DATA_OUT_31_port
                           , B2 => n5, ZN => n74);
   U33 : AOI22_X1 port map( A1 => DATA_IN(30), A2 => n6, B1 => DATA_OUT_30_port
                           , B2 => n5, ZN => n75);
   U32 : AOI22_X1 port map( A1 => DATA_IN(29), A2 => n6, B1 => DATA_OUT_29_port
                           , B2 => n5, ZN => n76);
   U30 : AOI22_X1 port map( A1 => DATA_IN(27), A2 => n6, B1 => DATA_OUT_27_port
                           , B2 => n5, ZN => n78);
   U29 : AOI22_X1 port map( A1 => DATA_IN(26), A2 => n6, B1 => DATA_OUT_26_port
                           , B2 => n5, ZN => n79);
   U28 : AOI22_X1 port map( A1 => DATA_IN(25), A2 => n6, B1 => DATA_OUT_25_port
                           , B2 => n5, ZN => n80);
   U27 : AOI22_X1 port map( A1 => DATA_IN(24), A2 => n6, B1 => DATA_OUT_24_port
                           , B2 => n5, ZN => n81);
   U26 : AOI22_X1 port map( A1 => DATA_IN(23), A2 => n6, B1 => DATA_OUT_23_port
                           , B2 => n4, ZN => n82);
   U25 : AOI22_X1 port map( A1 => DATA_IN(22), A2 => n6, B1 => DATA_OUT_22_port
                           , B2 => n4, ZN => n83);
   U24 : AOI22_X1 port map( A1 => DATA_IN(21), A2 => n6, B1 => DATA_OUT_21_port
                           , B2 => n4, ZN => n84);
   U23 : AOI22_X1 port map( A1 => DATA_IN(20), A2 => n6, B1 => DATA_OUT_20_port
                           , B2 => n4, ZN => n85);
   U21 : AOI22_X1 port map( A1 => DATA_IN(18), A2 => n7, B1 => DATA_OUT_18_port
                           , B2 => n4, ZN => n87);
   U20 : AOI22_X1 port map( A1 => DATA_IN(17), A2 => n7, B1 => DATA_OUT_17_port
                           , B2 => n4, ZN => n88);
   U19 : AOI22_X1 port map( A1 => DATA_IN(16), A2 => n7, B1 => DATA_OUT_16_port
                           , B2 => n4, ZN => n89);
   U18 : AOI22_X1 port map( A1 => DATA_IN(15), A2 => n7, B1 => DATA_OUT_15_port
                           , B2 => n4, ZN => n90);
   U17 : AOI22_X1 port map( A1 => DATA_IN(14), A2 => n7, B1 => DATA_OUT_14_port
                           , B2 => n4, ZN => n91);
   U16 : AOI22_X1 port map( A1 => DATA_IN(13), A2 => n7, B1 => DATA_OUT_13_port
                           , B2 => n4, ZN => n92);
   U15 : AOI22_X1 port map( A1 => DATA_IN(12), A2 => n7, B1 => DATA_OUT_12_port
                           , B2 => n4, ZN => n93);
   U14 : AOI22_X1 port map( A1 => DATA_IN(11), A2 => n7, B1 => DATA_OUT_11_port
                           , B2 => n3, ZN => n94);
   U13 : AOI22_X1 port map( A1 => DATA_IN(10), A2 => n7, B1 => DATA_OUT_10_port
                           , B2 => n3, ZN => n95);
   U12 : AOI22_X1 port map( A1 => DATA_IN(9), A2 => n7, B1 => DATA_OUT_9_port, 
                           B2 => n3, ZN => n96);
   U11 : AOI22_X1 port map( A1 => DATA_IN(8), A2 => n7, B1 => DATA_OUT_8_port, 
                           B2 => n3, ZN => n97);
   U35 : NOR2_X1 port map( A1 => n2, A2 => n5, ZN => n105);
   U36 : BUF_X1 port map( A => n105, Z => n7);
   U37 : BUF_X1 port map( A => n105, Z => n6);
   U38 : BUF_X1 port map( A => n105, Z => n8);
   U39 : BUF_X1 port map( A => n1, Z => n3);
   U40 : BUF_X1 port map( A => n1, Z => n4);
   U41 : BUF_X1 port map( A => n1, Z => n5);
   U42 : NOR2_X1 port map( A1 => EN, A2 => n2, ZN => n1);
   U43 : INV_X1 port map( A => RST, ZN => n2);
   U44 : INV_X1 port map( A => n106, ZN => n73);
   U45 : INV_X1 port map( A => n104, ZN => n72);
   U46 : INV_X1 port map( A => n103, ZN => n71);
   U47 : INV_X1 port map( A => n102, ZN => n70);
   U48 : INV_X1 port map( A => n101, ZN => n69);
   U49 : INV_X1 port map( A => n100, ZN => n68);
   U50 : INV_X1 port map( A => n99, ZN => n36);
   U51 : INV_X1 port map( A => n98, ZN => n33);
   U52 : INV_X1 port map( A => n97, ZN => n32);
   U53 : INV_X1 port map( A => n96, ZN => n31);
   U54 : INV_X1 port map( A => n95, ZN => n30);
   U55 : INV_X1 port map( A => n94, ZN => n29);
   U56 : INV_X1 port map( A => n93, ZN => n28);
   U57 : INV_X1 port map( A => n92, ZN => n27);
   U58 : INV_X1 port map( A => n91, ZN => n26);
   U59 : INV_X1 port map( A => n90, ZN => n25);
   U60 : INV_X1 port map( A => n89, ZN => n24);
   U61 : INV_X1 port map( A => n88, ZN => n23);
   U62 : INV_X1 port map( A => n87, ZN => n22);
   U63 : INV_X1 port map( A => n86, ZN => n21);
   U64 : INV_X1 port map( A => n85, ZN => n20);
   U65 : INV_X1 port map( A => n84, ZN => n19);
   U66 : INV_X1 port map( A => n83, ZN => n18);
   U67 : INV_X1 port map( A => n82, ZN => n17);
   U68 : INV_X1 port map( A => n81, ZN => n16);
   U69 : INV_X1 port map( A => n80, ZN => n15);
   U70 : INV_X1 port map( A => n79, ZN => n14);
   U71 : INV_X1 port map( A => n78, ZN => n13);
   U72 : INV_X1 port map( A => n77, ZN => n12);
   U73 : INV_X1 port map( A => n76, ZN => n11);
   U74 : INV_X1 port map( A => n75, ZN => n10);
   U75 : INV_X1 port map( A => n74, ZN => n9);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_2 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_2;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_2 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n_2219,
      n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, 
      n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, 
      n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, 
      n_2247, n_2248, n_2249, n_2250 : std_logic;

begin
   DATA_OUT <= ( n67, n65, n63, n61, n59, n57, n55, n53, n51, n49, n47, n45, 
      n43, n41, n39, n37, n35, n33, n31, n29, n27, n25, n23, n21, n19, n17, n15
      , n13, n11, n9, n7, n5 );
   
   U3 : BUF_X2 port map( A => n106, Z => n71);
   U4 : BUF_X2 port map( A => n106, Z => n72);
   U5 : BUF_X1 port map( A => n1, Z => n68);
   U6 : BUF_X1 port map( A => n1, Z => n69);
   U7 : BUF_X1 port map( A => n106, Z => n73);
   U8 : BUF_X1 port map( A => n1, Z => n70);
   U9 : AND2_X1 port map( A1 => n2, A2 => n74, ZN => n1);
   U10 : INV_X1 port map( A => n3, ZN => n2);
   U11 : INV_X1 port map( A => RST, ZN => n3);
   U44 : OR2_X1 port map( A1 => EN, A2 => n3, ZN => n74);
   U45 : INV_X1 port map( A => n74, ZN => n106);
   U46 : AOI22_X1 port map( A1 => n5, A2 => n71, B1 => DATA_IN(0), B2 => n68, 
                           ZN => n75);
   U47 : INV_X1 port map( A => n75, ZN => n139);
   U48 : AOI22_X1 port map( A1 => n7, A2 => n71, B1 => DATA_IN(1), B2 => n68, 
                           ZN => n76);
   U49 : INV_X1 port map( A => n76, ZN => n138);
   U50 : AOI22_X1 port map( A1 => n9, A2 => n71, B1 => DATA_IN(2), B2 => n68, 
                           ZN => n77);
   U51 : INV_X1 port map( A => n77, ZN => n137);
   U52 : AOI22_X1 port map( A1 => n11, A2 => n71, B1 => DATA_IN(3), B2 => n68, 
                           ZN => n78);
   U53 : INV_X1 port map( A => n78, ZN => n136);
   U54 : AOI22_X1 port map( A1 => n13, A2 => n71, B1 => DATA_IN(4), B2 => n68, 
                           ZN => n79);
   U55 : INV_X1 port map( A => n79, ZN => n135);
   U56 : AOI22_X1 port map( A1 => n15, A2 => n71, B1 => DATA_IN(5), B2 => n68, 
                           ZN => n80);
   U57 : INV_X1 port map( A => n80, ZN => n134);
   U58 : AOI22_X1 port map( A1 => n17, A2 => n71, B1 => DATA_IN(6), B2 => n68, 
                           ZN => n81);
   U59 : INV_X1 port map( A => n81, ZN => n133);
   U60 : AOI22_X1 port map( A1 => n19, A2 => n71, B1 => DATA_IN(7), B2 => n68, 
                           ZN => n82);
   U61 : INV_X1 port map( A => n82, ZN => n132);
   U62 : AOI22_X1 port map( A1 => n21, A2 => n71, B1 => DATA_IN(8), B2 => n68, 
                           ZN => n83);
   U63 : INV_X1 port map( A => n83, ZN => n131);
   U64 : AOI22_X1 port map( A1 => n23, A2 => n71, B1 => DATA_IN(9), B2 => n68, 
                           ZN => n84);
   U65 : INV_X1 port map( A => n84, ZN => n130);
   U66 : AOI22_X1 port map( A1 => n25, A2 => n71, B1 => DATA_IN(10), B2 => n68,
                           ZN => n85);
   U67 : INV_X1 port map( A => n85, ZN => n129);
   U68 : AOI22_X1 port map( A1 => n27, A2 => n71, B1 => DATA_IN(11), B2 => n68,
                           ZN => n86);
   U69 : INV_X1 port map( A => n86, ZN => n128);
   U70 : AOI22_X1 port map( A1 => n29, A2 => n72, B1 => DATA_IN(12), B2 => n69,
                           ZN => n87);
   U71 : INV_X1 port map( A => n87, ZN => n127);
   U72 : AOI22_X1 port map( A1 => n31, A2 => n72, B1 => DATA_IN(13), B2 => n69,
                           ZN => n88);
   U73 : INV_X1 port map( A => n88, ZN => n126);
   U74 : AOI22_X1 port map( A1 => n33, A2 => n72, B1 => DATA_IN(14), B2 => n69,
                           ZN => n89);
   U75 : INV_X1 port map( A => n89, ZN => n125);
   U76 : AOI22_X1 port map( A1 => n35, A2 => n72, B1 => DATA_IN(15), B2 => n69,
                           ZN => n90);
   U77 : INV_X1 port map( A => n90, ZN => n124);
   U78 : AOI22_X1 port map( A1 => n37, A2 => n72, B1 => DATA_IN(16), B2 => n69,
                           ZN => n91);
   U79 : INV_X1 port map( A => n91, ZN => n123);
   U80 : AOI22_X1 port map( A1 => n39, A2 => n72, B1 => DATA_IN(17), B2 => n69,
                           ZN => n92);
   U81 : INV_X1 port map( A => n92, ZN => n122);
   U82 : AOI22_X1 port map( A1 => n41, A2 => n72, B1 => DATA_IN(18), B2 => n69,
                           ZN => n93);
   U83 : INV_X1 port map( A => n93, ZN => n121);
   U84 : AOI22_X1 port map( A1 => n43, A2 => n72, B1 => DATA_IN(19), B2 => n69,
                           ZN => n94);
   U85 : INV_X1 port map( A => n94, ZN => n120);
   U86 : AOI22_X1 port map( A1 => n45, A2 => n72, B1 => DATA_IN(20), B2 => n69,
                           ZN => n95);
   U87 : INV_X1 port map( A => n95, ZN => n119);
   U88 : AOI22_X1 port map( A1 => n47, A2 => n72, B1 => DATA_IN(21), B2 => n69,
                           ZN => n96);
   U89 : INV_X1 port map( A => n96, ZN => n118);
   U90 : AOI22_X1 port map( A1 => n49, A2 => n72, B1 => DATA_IN(22), B2 => n69,
                           ZN => n97);
   U91 : INV_X1 port map( A => n97, ZN => n117);
   U92 : AOI22_X1 port map( A1 => n51, A2 => n72, B1 => DATA_IN(23), B2 => n69,
                           ZN => n98);
   U93 : INV_X1 port map( A => n98, ZN => n116);
   U94 : AOI22_X1 port map( A1 => n53, A2 => n73, B1 => DATA_IN(24), B2 => n70,
                           ZN => n99);
   U95 : INV_X1 port map( A => n99, ZN => n115);
   U96 : AOI22_X1 port map( A1 => n55, A2 => n73, B1 => DATA_IN(25), B2 => n70,
                           ZN => n100);
   U97 : INV_X1 port map( A => n100, ZN => n114);
   U98 : AOI22_X1 port map( A1 => n57, A2 => n73, B1 => DATA_IN(26), B2 => n70,
                           ZN => n101);
   U99 : INV_X1 port map( A => n101, ZN => n113);
   U100 : AOI22_X1 port map( A1 => n59, A2 => n73, B1 => DATA_IN(27), B2 => n70
                           , ZN => n102);
   U101 : INV_X1 port map( A => n102, ZN => n112);
   U102 : AOI22_X1 port map( A1 => n61, A2 => n73, B1 => DATA_IN(28), B2 => n70
                           , ZN => n103);
   U103 : INV_X1 port map( A => n103, ZN => n111);
   U104 : AOI22_X1 port map( A1 => n63, A2 => n73, B1 => DATA_IN(29), B2 => n70
                           , ZN => n104);
   U105 : INV_X1 port map( A => n104, ZN => n110);
   U106 : AOI22_X1 port map( A1 => n65, A2 => n73, B1 => DATA_IN(30), B2 => n70
                           , ZN => n105);
   U107 : INV_X1 port map( A => n105, ZN => n109);
   U108 : AOI22_X1 port map( A1 => n67, A2 => n73, B1 => DATA_IN(31), B2 => n70
                           , ZN => n107);
   U109 : INV_X1 port map( A => n107, ZN => n108);
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n108, CK => CLK, Q => n67, QN 
                           => n_2219);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n109, CK => CLK, Q => n65, QN 
                           => n_2220);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n110, CK => CLK, Q => n63, QN 
                           => n_2221);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n111, CK => CLK, Q => n61, QN 
                           => n_2222);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n112, CK => CLK, Q => n59, QN 
                           => n_2223);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n113, CK => CLK, Q => n57, QN 
                           => n_2224);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n114, CK => CLK, Q => n55, QN 
                           => n_2225);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n115, CK => CLK, Q => n53, QN 
                           => n_2226);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n116, CK => CLK, Q => n51, QN 
                           => n_2227);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n117, CK => CLK, Q => n49, QN 
                           => n_2228);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n118, CK => CLK, Q => n47, QN 
                           => n_2229);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n119, CK => CLK, Q => n45, QN 
                           => n_2230);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n120, CK => CLK, Q => n43, QN 
                           => n_2231);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n121, CK => CLK, Q => n41, QN 
                           => n_2232);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n122, CK => CLK, Q => n39, QN 
                           => n_2233);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n123, CK => CLK, Q => n37, QN 
                           => n_2234);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n124, CK => CLK, Q => n35, QN 
                           => n_2235);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n125, CK => CLK, Q => n33, QN 
                           => n_2236);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n126, CK => CLK, Q => n31, QN 
                           => n_2237);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n127, CK => CLK, Q => n29, QN 
                           => n_2238);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n128, CK => CLK, Q => n27, QN 
                           => n_2239);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n129, CK => CLK, Q => n25, QN 
                           => n_2240);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n130, CK => CLK, Q => n23, QN =>
                           n_2241);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n131, CK => CLK, Q => n21, QN =>
                           n_2242);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n132, CK => CLK, Q => n19, QN =>
                           n_2243);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n133, CK => CLK, Q => n17, QN =>
                           n_2244);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n134, CK => CLK, Q => n15, QN =>
                           n_2245);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n135, CK => CLK, Q => n13, QN =>
                           n_2246);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n136, CK => CLK, Q => n11, QN =>
                           n_2247);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n137, CK => CLK, Q => n9, QN => 
                           n_2248);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n138, CK => CLK, Q => n7, QN => 
                           n_2249);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n139, CK => CLK, Q => n5, QN => 
                           n_2250);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_3 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_3;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_3 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, net51629, net51627, 
      net51625, net51635, net51633, net51631, n1, n2, n3, n4, n5, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n73, n75, n77, n79, n81, n83, n84, n85, n86, n87, n88
      , n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102
      , n103, n104, n105, n106, n107, n108, n109, n_2251, n_2252, n_2253, 
      n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, 
      n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, 
      n_2272, n_2273, n_2274, n_2275, n_2276, n_2277 : std_logic;

begin
   DATA_OUT <= ( DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, n83, n81, n79, n77, 
      n75, n73 );
   
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n98, CK => CLK, Q => 
                           DATA_OUT_30_port, QN => n_2251);
   DATA_OUT_reg_20_inst : DFF_X2 port map( D => n102, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_2252);
   DATA_OUT_reg_23_inst : DFF_X2 port map( D => n60, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_2253);
   DATA_OUT_reg_17_inst : DFF_X2 port map( D => n57, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_2254);
   DATA_OUT_reg_19_inst : DFF_X2 port map( D => n54, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_2255);
   DATA_OUT_reg_18_inst : DFF_X2 port map( D => n51, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_2256);
   DATA_OUT_reg_8_inst : DFF_X2 port map( D => n42, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n_2257);
   DATA_OUT_reg_6_inst : DFF_X2 port map( D => n48, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n_2258);
   DATA_OUT_reg_27_inst : DFF_X2 port map( D => n99, CK => CLK, Q => 
                           DATA_OUT_27_port, QN => n_2259);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n100, CK => CLK, Q => 
                           DATA_OUT_26_port, QN => n_2260);
   DATA_OUT_reg_11_inst : DFF_X2 port map( D => n106, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n_2261);
   DATA_OUT_reg_7_inst : DFF_X2 port map( D => n39, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n_2262);
   DATA_OUT_reg_28_inst : DFF_X2 port map( D => n45, CK => CLK, Q => 
                           DATA_OUT_28_port, QN => n_2263);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n103, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n_2264);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n101, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_2265);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n104, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n_2266);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n105, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n_2267);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n107, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n_2268);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n108, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n_2269);
   U3 : OR2_X1 port map( A1 => n1, A2 => n24, ZN => n14);
   U4 : BUF_X1 port map( A => n71, Z => net51631);
   U5 : AND2_X2 port map( A1 => n69, A2 => n68, ZN => n71);
   U6 : INV_X1 port map( A => n10, ZN => n11);
   U8 : NAND2_X1 port map( A1 => DATA_OUT_29_port, A2 => net51629, ZN => n7);
   U9 : NAND2_X1 port map( A1 => DATA_IN(29), A2 => net51635, ZN => n8);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n9);
   U11 : INV_X1 port map( A => n71, ZN => n10);
   U12 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => n12);
   U13 : NAND2_X1 port map( A1 => DATA_IN(15), A2 => n11, ZN => n13);
   U14 : CLKBUF_X3 port map( A => n67, Z => net51625);
   U15 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n15);
   U16 : NAND2_X1 port map( A1 => DATA_IN(21), A2 => n11, ZN => n16);
   U17 : OR2_X4 port map( A1 => n2, A2 => n24, ZN => n17);
   U18 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => n18);
   U19 : NAND2_X1 port map( A1 => DATA_IN(22), A2 => net51633, ZN => n19);
   U20 : OR2_X4 port map( A1 => n3, A2 => n24, ZN => n20);
   U21 : BUF_X1 port map( A => n71, Z => net51633);
   U22 : NAND2_X1 port map( A1 => n75, A2 => net51625, ZN => n21);
   U23 : NAND2_X1 port map( A1 => DATA_IN(1), A2 => net51631, ZN => n22);
   U24 : NAND2_X1 port map( A1 => n22, A2 => n21, ZN => n23);
   U25 : CLKBUF_X1 port map( A => n71, Z => net51635);
   U26 : INV_X1 port map( A => n67, ZN => n24);
   U27 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => n25);
   U28 : NAND2_X1 port map( A1 => DATA_IN(16), A2 => n11, ZN => n26);
   U29 : OR2_X4 port map( A1 => n4, A2 => n24, ZN => n27);
   U30 : NAND2_X1 port map( A1 => n79, A2 => net51625, ZN => n28);
   U31 : NAND2_X1 port map( A1 => DATA_IN(3), A2 => net51631, ZN => n29);
   U32 : NAND2_X1 port map( A1 => n29, A2 => n28, ZN => n30);
   U33 : NAND2_X1 port map( A1 => n77, A2 => net51625, ZN => n31);
   U34 : NAND2_X1 port map( A1 => DATA_IN(2), A2 => net51631, ZN => n32);
   U35 : NAND2_X1 port map( A1 => n32, A2 => n31, ZN => n33);
   U36 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => n34);
   U37 : NAND2_X1 port map( A1 => DATA_IN(24), A2 => n11, ZN => n35);
   U38 : OR2_X4 port map( A1 => n5, A2 => n24, ZN => n36);
   U39 : NAND2_X1 port map( A1 => DATA_OUT_7_port, A2 => net51625, ZN => n37);
   U40 : NAND2_X1 port map( A1 => DATA_IN(7), A2 => net51631, ZN => n38);
   U41 : NAND2_X1 port map( A1 => n38, A2 => n37, ZN => n39);
   U42 : NAND2_X1 port map( A1 => DATA_OUT_8_port, A2 => net51625, ZN => n40);
   U43 : NAND2_X1 port map( A1 => DATA_IN(8), A2 => net51631, ZN => n41);
   U44 : NAND2_X1 port map( A1 => n41, A2 => n40, ZN => n42);
   U45 : NAND2_X1 port map( A1 => DATA_OUT_28_port, A2 => net51629, ZN => n43);
   U46 : NAND2_X1 port map( A1 => DATA_IN(28), A2 => net51635, ZN => n44);
   U47 : NAND2_X1 port map( A1 => n44, A2 => n43, ZN => n45);
   U48 : NAND2_X1 port map( A1 => DATA_OUT_6_port, A2 => net51625, ZN => n46);
   U49 : NAND2_X1 port map( A1 => DATA_IN(6), A2 => net51631, ZN => n47);
   U50 : NAND2_X1 port map( A1 => n47, A2 => n46, ZN => n48);
   U51 : NAND2_X1 port map( A1 => DATA_OUT_18_port, A2 => net51627, ZN => n49);
   U52 : NAND2_X1 port map( A1 => DATA_IN(18), A2 => net51633, ZN => n50);
   U53 : NAND2_X1 port map( A1 => n50, A2 => n49, ZN => n51);
   U54 : NAND2_X1 port map( A1 => DATA_OUT_19_port, A2 => net51627, ZN => n52);
   U55 : NAND2_X1 port map( A1 => DATA_IN(19), A2 => net51633, ZN => n53);
   U56 : NAND2_X1 port map( A1 => n53, A2 => n52, ZN => n54);
   U57 : NAND2_X1 port map( A1 => DATA_OUT_17_port, A2 => net51627, ZN => n55);
   U58 : NAND2_X1 port map( A1 => DATA_IN(17), A2 => net51633, ZN => n56);
   U59 : NAND2_X1 port map( A1 => n56, A2 => n55, ZN => n57);
   U60 : NAND2_X1 port map( A1 => DATA_OUT_23_port, A2 => net51627, ZN => n58);
   U61 : NAND2_X1 port map( A1 => DATA_IN(23), A2 => net51633, ZN => n59);
   U62 : NAND2_X1 port map( A1 => n59, A2 => n58, ZN => n60);
   U63 : NAND2_X1 port map( A1 => n73, A2 => net51625, ZN => n61);
   U64 : NAND2_X1 port map( A1 => DATA_IN(0), A2 => net51631, ZN => n62);
   U65 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => n63);
   U66 : NAND2_X1 port map( A1 => n83, A2 => net51625, ZN => n64);
   U67 : NAND2_X1 port map( A1 => DATA_IN(5), A2 => net51631, ZN => n65);
   U68 : NAND2_X1 port map( A1 => n65, A2 => n64, ZN => n66);
   U69 : AOI22_X1 port map( A1 => DATA_IN(20), A2 => n71, B1 => net51627, B2 =>
                           DATA_OUT_20_port, ZN => n91);
   U70 : BUF_X2 port map( A => n67, Z => net51629);
   U71 : AOI22_X1 port map( A1 => DATA_IN(4), A2 => n71, B1 => n81, B2 => n67, 
                           ZN => n84);
   U72 : INV_X2 port map( A => n68, ZN => n67);
   U73 : AOI22_X1 port map( A1 => DATA_IN(30), A2 => n71, B1 => net51629, B2 =>
                           DATA_OUT_30_port, ZN => n95);
   U74 : AOI22_X1 port map( A1 => DATA_IN(14), A2 => n71, B1 => net51627, B2 =>
                           DATA_OUT_14_port, ZN => n90);
   U75 : BUF_X2 port map( A => n67, Z => net51627);
   U76 : AOI22_X1 port map( A1 => DATA_IN(27), A2 => n71, B1 => net51629, B2 =>
                           DATA_OUT_27_port, ZN => n94);
   U77 : AOI22_X1 port map( A1 => DATA_IN(9), A2 => n71, B1 => net51625, B2 => 
                           DATA_OUT_9_port, ZN => n85);
   U78 : AOI22_X1 port map( A1 => DATA_IN(12), A2 => n71, B1 => n67, B2 => 
                           DATA_OUT_12_port, ZN => n88);
   U79 : AOI22_X1 port map( A1 => DATA_IN(26), A2 => n71, B1 => net51629, B2 =>
                           DATA_OUT_26_port, ZN => n93);
   U80 : AOI22_X1 port map( A1 => DATA_IN(10), A2 => n71, B1 => net51625, B2 =>
                           DATA_OUT_10_port, ZN => n86);
   U81 : AOI22_X1 port map( A1 => DATA_IN(13), A2 => n71, B1 => n67, B2 => 
                           DATA_OUT_13_port, ZN => n89);
   U82 : AOI22_X1 port map( A1 => DATA_IN(25), A2 => n71, B1 => net51629, B2 =>
                           DATA_OUT_25_port, ZN => n92);
   U83 : AOI22_X1 port map( A1 => DATA_IN(11), A2 => n71, B1 => n67, B2 => 
                           DATA_OUT_11_port, ZN => n87);
   U84 : INV_X1 port map( A => n70, ZN => n69);
   U85 : INV_X1 port map( A => RST, ZN => n70);
   U86 : OR2_X1 port map( A1 => EN, A2 => n70, ZN => n68);
   U93 : INV_X1 port map( A => n84, ZN => n109);
   U94 : INV_X1 port map( A => n85, ZN => n108);
   U95 : INV_X1 port map( A => n86, ZN => n107);
   U96 : INV_X1 port map( A => n87, ZN => n106);
   U97 : INV_X1 port map( A => n88, ZN => n105);
   U98 : INV_X1 port map( A => n89, ZN => n104);
   U99 : INV_X1 port map( A => n90, ZN => n103);
   U100 : INV_X1 port map( A => n91, ZN => n102);
   U101 : INV_X1 port map( A => n92, ZN => n101);
   U102 : INV_X1 port map( A => n93, ZN => n100);
   U103 : INV_X1 port map( A => n94, ZN => n99);
   U104 : INV_X1 port map( A => n95, ZN => n98);
   U105 : AOI22_X1 port map( A1 => DATA_OUT_31_port, A2 => net51629, B1 => 
                           DATA_IN(31), B2 => net51635, ZN => n96);
   U106 : INV_X1 port map( A => n96, ZN => n97);
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n97, CK => CLK, Q => 
                           DATA_OUT_31_port, QN => n_2270);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n63, CK => CLK, Q => n73, QN => 
                           n_2271);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n23, CK => CLK, Q => n75, QN => 
                           n_2272);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n30, CK => CLK, Q => n79, QN => 
                           n_2273);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n33, CK => CLK, Q => n77, QN => 
                           n_2274);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n66, CK => CLK, Q => n83, QN => 
                           n_2275);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n25, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n4);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n12, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n1);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n15, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n2);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n18, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n3);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n34, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n5);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n109, CK => CLK, Q => n81, QN =>
                           n_2276);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n9, CK => CLK, Q => 
                           DATA_OUT_29_port, QN => n_2277);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT5_2 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 downto 
         0);  DATA_OUT : out std_logic_vector (4 downto 0));

end REG_GENERIC_NBIT5_2;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT5_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n_2278, n_2279, n_2280, n_2281, n_2282 : std_logic;

begin
   DATA_OUT <= ( DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, 
      DATA_OUT_1_port, DATA_OUT_0_port );
   
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n11, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_2278);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n12, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_2279);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n13, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_2280);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n14, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_2281);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n15, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_2282);
   U3 : AND2_X1 port map( A1 => n2, A2 => n4, ZN => n1);
   U4 : INV_X1 port map( A => n3, ZN => n2);
   U5 : INV_X1 port map( A => RST, ZN => n3);
   U6 : OR2_X1 port map( A1 => EN, A2 => n3, ZN => n4);
   U7 : INV_X1 port map( A => n4, ZN => n9);
   U8 : AOI22_X1 port map( A1 => DATA_OUT_0_port, A2 => n9, B1 => DATA_IN(0), 
                           B2 => n1, ZN => n5);
   U9 : INV_X1 port map( A => n5, ZN => n15);
   U10 : AOI22_X1 port map( A1 => DATA_OUT_1_port, A2 => n9, B1 => DATA_IN(1), 
                           B2 => n1, ZN => n6);
   U11 : INV_X1 port map( A => n6, ZN => n14);
   U12 : AOI22_X1 port map( A1 => DATA_OUT_2_port, A2 => n9, B1 => DATA_IN(2), 
                           B2 => n1, ZN => n7);
   U13 : INV_X1 port map( A => n7, ZN => n13);
   U14 : AOI22_X1 port map( A1 => DATA_OUT_3_port, A2 => n9, B1 => DATA_IN(3), 
                           B2 => n1, ZN => n8);
   U15 : INV_X1 port map( A => n8, ZN => n12);
   U16 : AOI22_X1 port map( A1 => DATA_OUT_4_port, A2 => n9, B1 => DATA_IN(4), 
                           B2 => n1, ZN => n10);
   U17 : INV_X1 port map( A => n10, ZN => n11);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT5_0 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 downto 
         0);  DATA_OUT : out std_logic_vector (4 downto 0));

end REG_GENERIC_NBIT5_0;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n9, n14, n15, n16, n17, n18, n19
      , n_2283, n_2284, n_2285, n_2286, n_2287 : std_logic;

begin
   DATA_OUT <= ( DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, 
      DATA_OUT_1_port, DATA_OUT_0_port );
   
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n3, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_2283);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n4, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_2284);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n5, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_2285);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n6, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_2286);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n9, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_2287);
   U7 : AOI22_X1 port map( A1 => DATA_IN(4), A2 => n18, B1 => DATA_OUT_4_port, 
                           B2 => n1, ZN => n14);
   U6 : AOI22_X1 port map( A1 => DATA_IN(3), A2 => n18, B1 => DATA_OUT_3_port, 
                           B2 => n1, ZN => n15);
   U5 : AOI22_X1 port map( A1 => DATA_IN(2), A2 => n18, B1 => DATA_OUT_2_port, 
                           B2 => n1, ZN => n16);
   U4 : AOI22_X1 port map( A1 => DATA_IN(1), A2 => n18, B1 => DATA_OUT_1_port, 
                           B2 => n1, ZN => n17);
   U3 : AOI22_X1 port map( A1 => DATA_IN(0), A2 => n18, B1 => DATA_OUT_0_port, 
                           B2 => n1, ZN => n19);
   U8 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => n18);
   U9 : NOR2_X1 port map( A1 => EN, A2 => n2, ZN => n1);
   U10 : INV_X1 port map( A => RST, ZN => n2);
   U11 : INV_X1 port map( A => n19, ZN => n9);
   U12 : INV_X1 port map( A => n17, ZN => n6);
   U13 : INV_X1 port map( A => n16, ZN => n5);
   U14 : INV_X1 port map( A => n15, ZN => n4);
   U15 : INV_X1 port map( A => n14, ZN => n3);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT26 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (25 downto
         0);  DATA_OUT : out std_logic_vector (25 downto 0));

end REG_GENERIC_NBIT26;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_25_port, DATA_OUT_24_port, DATA_OUT_23_port, 
      DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, DATA_OUT_19_port, 
      DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, DATA_OUT_15_port, 
      DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, DATA_OUT_11_port, 
      DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, DATA_OUT_7_port, 
      DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, DATA_OUT_3_port, 
      DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port, n1, n2, n3, n4, n5, n6
      , n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n_2288, 
      n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, 
      n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, 
      n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313 : std_logic;

begin
   DATA_OUT <= ( DATA_OUT_25_port, DATA_OUT_24_port, DATA_OUT_23_port, 
      DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, DATA_OUT_19_port, 
      DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, DATA_OUT_15_port, 
      DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, DATA_OUT_11_port, 
      DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, DATA_OUT_7_port, 
      DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, DATA_OUT_3_port, 
      DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port );
   
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n38, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_2288);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n39, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n_2289);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n40, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_2290);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n41, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n_2291);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n42, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n_2292);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n43, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_2293);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n44, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_2294);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n45, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_2295);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n46, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_2296);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n47, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n_2297);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n48, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n_2298);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n49, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n_2299);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n50, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n_2300);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n51, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n_2301);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n52, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n_2302);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n53, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n_2303);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n54, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n_2304);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n55, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n_2305);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n56, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n_2306);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n57, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n_2307);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n58, CK => CLK, Q => 
                           DATA_OUT_5_port, QN => n_2308);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n59, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_2309);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n60, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_2310);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n61, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_2311);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n62, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_2312);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n63, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_2313);
   U3 : CLKBUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X2 port map( A => n36, Z => n7);
   U5 : BUF_X2 port map( A => n36, Z => n8);
   U6 : BUF_X1 port map( A => n1, Z => n5);
   U7 : BUF_X1 port map( A => n1, Z => n4);
   U8 : CLKBUF_X1 port map( A => n36, Z => n9);
   U9 : AND2_X1 port map( A1 => n2, A2 => n10, ZN => n1);
   U10 : INV_X1 port map( A => n3, ZN => n2);
   U11 : INV_X1 port map( A => RST, ZN => n3);
   U12 : OR2_X1 port map( A1 => EN, A2 => n3, ZN => n10);
   U13 : INV_X1 port map( A => n10, ZN => n36);
   U14 : AOI22_X1 port map( A1 => DATA_OUT_0_port, A2 => n7, B1 => DATA_IN(0), 
                           B2 => n6, ZN => n11);
   U15 : INV_X1 port map( A => n11, ZN => n63);
   U16 : AOI22_X1 port map( A1 => DATA_OUT_1_port, A2 => n7, B1 => DATA_IN(1), 
                           B2 => n6, ZN => n12);
   U17 : INV_X1 port map( A => n12, ZN => n62);
   U18 : AOI22_X1 port map( A1 => DATA_OUT_2_port, A2 => n7, B1 => DATA_IN(2), 
                           B2 => n5, ZN => n13);
   U19 : INV_X1 port map( A => n13, ZN => n61);
   U20 : AOI22_X1 port map( A1 => DATA_OUT_3_port, A2 => n7, B1 => DATA_IN(3), 
                           B2 => n5, ZN => n14);
   U21 : INV_X1 port map( A => n14, ZN => n60);
   U22 : AOI22_X1 port map( A1 => DATA_OUT_4_port, A2 => n7, B1 => DATA_IN(4), 
                           B2 => n5, ZN => n15);
   U23 : INV_X1 port map( A => n15, ZN => n59);
   U24 : AOI22_X1 port map( A1 => DATA_OUT_5_port, A2 => n7, B1 => DATA_IN(5), 
                           B2 => n5, ZN => n16);
   U25 : INV_X1 port map( A => n16, ZN => n58);
   U26 : AOI22_X1 port map( A1 => DATA_OUT_6_port, A2 => n7, B1 => DATA_IN(6), 
                           B2 => n5, ZN => n17);
   U27 : INV_X1 port map( A => n17, ZN => n57);
   U28 : AOI22_X1 port map( A1 => DATA_OUT_7_port, A2 => n7, B1 => DATA_IN(7), 
                           B2 => n5, ZN => n18);
   U29 : INV_X1 port map( A => n18, ZN => n56);
   U30 : AOI22_X1 port map( A1 => DATA_OUT_8_port, A2 => n7, B1 => DATA_IN(8), 
                           B2 => n5, ZN => n19);
   U31 : INV_X1 port map( A => n19, ZN => n55);
   U32 : AOI22_X1 port map( A1 => DATA_OUT_9_port, A2 => n7, B1 => DATA_IN(9), 
                           B2 => n5, ZN => n20);
   U33 : INV_X1 port map( A => n20, ZN => n54);
   U34 : AOI22_X1 port map( A1 => DATA_OUT_10_port, A2 => n7, B1 => DATA_IN(10)
                           , B2 => n5, ZN => n21);
   U35 : INV_X1 port map( A => n21, ZN => n53);
   U36 : AOI22_X1 port map( A1 => DATA_OUT_11_port, A2 => n7, B1 => DATA_IN(11)
                           , B2 => n5, ZN => n22);
   U37 : INV_X1 port map( A => n22, ZN => n52);
   U38 : AOI22_X1 port map( A1 => DATA_OUT_12_port, A2 => n8, B1 => DATA_IN(12)
                           , B2 => n5, ZN => n23);
   U39 : INV_X1 port map( A => n23, ZN => n51);
   U40 : AOI22_X1 port map( A1 => DATA_OUT_13_port, A2 => n8, B1 => DATA_IN(13)
                           , B2 => n5, ZN => n24);
   U41 : INV_X1 port map( A => n24, ZN => n50);
   U42 : AOI22_X1 port map( A1 => DATA_OUT_14_port, A2 => n8, B1 => DATA_IN(14)
                           , B2 => n4, ZN => n25);
   U43 : INV_X1 port map( A => n25, ZN => n49);
   U44 : AOI22_X1 port map( A1 => DATA_OUT_15_port, A2 => n8, B1 => DATA_IN(15)
                           , B2 => n4, ZN => n26);
   U45 : INV_X1 port map( A => n26, ZN => n48);
   U46 : AOI22_X1 port map( A1 => DATA_OUT_16_port, A2 => n8, B1 => DATA_IN(16)
                           , B2 => n4, ZN => n27);
   U47 : INV_X1 port map( A => n27, ZN => n47);
   U48 : AOI22_X1 port map( A1 => DATA_OUT_17_port, A2 => n8, B1 => DATA_IN(17)
                           , B2 => n4, ZN => n28);
   U49 : INV_X1 port map( A => n28, ZN => n46);
   U50 : AOI22_X1 port map( A1 => DATA_OUT_18_port, A2 => n8, B1 => DATA_IN(18)
                           , B2 => n4, ZN => n29);
   U51 : INV_X1 port map( A => n29, ZN => n45);
   U52 : AOI22_X1 port map( A1 => DATA_OUT_19_port, A2 => n8, B1 => DATA_IN(19)
                           , B2 => n4, ZN => n30);
   U53 : INV_X1 port map( A => n30, ZN => n44);
   U54 : AOI22_X1 port map( A1 => DATA_OUT_20_port, A2 => n8, B1 => DATA_IN(20)
                           , B2 => n4, ZN => n31);
   U55 : INV_X1 port map( A => n31, ZN => n43);
   U56 : AOI22_X1 port map( A1 => DATA_OUT_21_port, A2 => n8, B1 => DATA_IN(21)
                           , B2 => n4, ZN => n32);
   U57 : INV_X1 port map( A => n32, ZN => n42);
   U58 : AOI22_X1 port map( A1 => DATA_OUT_22_port, A2 => n8, B1 => DATA_IN(22)
                           , B2 => n4, ZN => n33);
   U59 : INV_X1 port map( A => n33, ZN => n41);
   U60 : AOI22_X1 port map( A1 => DATA_OUT_23_port, A2 => n8, B1 => DATA_IN(23)
                           , B2 => n4, ZN => n34);
   U61 : INV_X1 port map( A => n34, ZN => n40);
   U62 : AOI22_X1 port map( A1 => DATA_OUT_24_port, A2 => n9, B1 => DATA_IN(24)
                           , B2 => n4, ZN => n35);
   U63 : INV_X1 port map( A => n35, ZN => n39);
   U64 : AOI22_X1 port map( A1 => DATA_OUT_25_port, A2 => n9, B1 => DATA_IN(25)
                           , B2 => n4, ZN => n37);
   U65 : INV_X1 port map( A => n37, ZN => n38);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_5 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_5;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n35, n36, n38, n68, n69, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88
      , n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102
      , n103, n104, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, 
      n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, 
      n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, 
      n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345 : std_logic;

begin
   DATA_OUT <= ( DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port );
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n11, CK => CLK, Q => 
                           DATA_OUT_31_port, QN => n_2314);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n12, CK => CLK, Q => 
                           DATA_OUT_30_port, QN => n_2315);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n13, CK => CLK, Q => 
                           DATA_OUT_29_port, QN => n_2316);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n14, CK => CLK, Q => 
                           DATA_OUT_28_port, QN => n_2317);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n15, CK => CLK, Q => 
                           DATA_OUT_27_port, QN => n_2318);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n16, CK => CLK, Q => 
                           DATA_OUT_26_port, QN => n_2319);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n17, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_2320);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n18, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n_2321);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n19, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_2322);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n20, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n_2323);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n21, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n_2324);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n22, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_2325);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n23, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_2326);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n24, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_2327);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n25, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_2328);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n26, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n_2329);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n27, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n_2330);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n28, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n_2331);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n29, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n_2332);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n30, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n_2333);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n31, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n_2334);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n32, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n_2335);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n33, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n_2336);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n35, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n_2337);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n36, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n_2338);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n38, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n_2339);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT_5_port, QN => n_2340);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_2341);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_2342);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_2343);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_2344);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_2345);
   U10 : AOI22_X1 port map( A1 => DATA_IN(7), A2 => n5, B1 => DATA_OUT_7_port, 
                           B2 => n8, ZN => n98);
   U9 : AOI22_X1 port map( A1 => DATA_IN(6), A2 => n5, B1 => DATA_OUT_6_port, 
                           B2 => n8, ZN => n99);
   U8 : AOI22_X1 port map( A1 => DATA_IN(5), A2 => n5, B1 => DATA_OUT_5_port, 
                           B2 => n8, ZN => n100);
   U7 : AOI22_X1 port map( A1 => DATA_IN(4), A2 => n5, B1 => DATA_OUT_4_port, 
                           B2 => n8, ZN => n101);
   U6 : AOI22_X1 port map( A1 => DATA_IN(3), A2 => n5, B1 => DATA_OUT_3_port, 
                           B2 => n8, ZN => n102);
   U4 : AOI22_X1 port map( A1 => DATA_IN(1), A2 => n5, B1 => DATA_OUT_1_port, 
                           B2 => n8, ZN => n103);
   U3 : AOI22_X1 port map( A1 => DATA_IN(0), A2 => n5, B1 => DATA_OUT_0_port, 
                           B2 => n8, ZN => n104);
   U34 : AOI22_X1 port map( A1 => DATA_IN(31), A2 => n3, B1 => DATA_OUT_31_port
                           , B2 => n6, ZN => n74);
   U33 : AOI22_X1 port map( A1 => DATA_IN(30), A2 => n3, B1 => DATA_OUT_30_port
                           , B2 => n6, ZN => n75);
   U32 : AOI22_X1 port map( A1 => DATA_IN(29), A2 => n3, B1 => DATA_OUT_29_port
                           , B2 => n6, ZN => n76);
   U31 : AOI22_X1 port map( A1 => DATA_IN(28), A2 => n3, B1 => DATA_OUT_28_port
                           , B2 => n6, ZN => n77);
   U30 : AOI22_X1 port map( A1 => DATA_IN(27), A2 => n3, B1 => DATA_OUT_27_port
                           , B2 => n6, ZN => n78);
   U29 : AOI22_X1 port map( A1 => DATA_IN(26), A2 => n3, B1 => DATA_OUT_26_port
                           , B2 => n6, ZN => n79);
   U28 : AOI22_X1 port map( A1 => DATA_IN(25), A2 => n3, B1 => DATA_OUT_25_port
                           , B2 => n6, ZN => n80);
   U27 : AOI22_X1 port map( A1 => DATA_IN(24), A2 => n3, B1 => DATA_OUT_24_port
                           , B2 => n6, ZN => n81);
   U26 : AOI22_X1 port map( A1 => DATA_IN(23), A2 => n3, B1 => DATA_OUT_23_port
                           , B2 => n6, ZN => n82);
   U25 : AOI22_X1 port map( A1 => DATA_IN(22), A2 => n3, B1 => DATA_OUT_22_port
                           , B2 => n6, ZN => n83);
   U24 : AOI22_X1 port map( A1 => DATA_IN(21), A2 => n3, B1 => DATA_OUT_21_port
                           , B2 => n6, ZN => n84);
   U23 : AOI22_X1 port map( A1 => DATA_IN(20), A2 => n3, B1 => DATA_OUT_20_port
                           , B2 => n6, ZN => n85);
   U22 : AOI22_X1 port map( A1 => DATA_IN(19), A2 => n4, B1 => DATA_OUT_19_port
                           , B2 => n7, ZN => n86);
   U21 : AOI22_X1 port map( A1 => DATA_IN(18), A2 => n4, B1 => DATA_OUT_18_port
                           , B2 => n7, ZN => n87);
   U20 : AOI22_X1 port map( A1 => DATA_IN(17), A2 => n4, B1 => DATA_OUT_17_port
                           , B2 => n7, ZN => n88);
   U19 : AOI22_X1 port map( A1 => DATA_IN(16), A2 => n4, B1 => DATA_OUT_16_port
                           , B2 => n7, ZN => n89);
   U18 : AOI22_X1 port map( A1 => DATA_IN(15), A2 => n4, B1 => DATA_OUT_15_port
                           , B2 => n7, ZN => n90);
   U17 : AOI22_X1 port map( A1 => DATA_IN(14), A2 => n4, B1 => DATA_OUT_14_port
                           , B2 => n7, ZN => n91);
   U16 : AOI22_X1 port map( A1 => DATA_IN(13), A2 => n4, B1 => DATA_OUT_13_port
                           , B2 => n7, ZN => n92);
   U15 : AOI22_X1 port map( A1 => DATA_IN(12), A2 => n4, B1 => DATA_OUT_12_port
                           , B2 => n7, ZN => n93);
   U14 : AOI22_X1 port map( A1 => DATA_IN(11), A2 => n4, B1 => DATA_OUT_11_port
                           , B2 => n7, ZN => n94);
   U13 : AOI22_X1 port map( A1 => DATA_IN(10), A2 => n4, B1 => DATA_OUT_10_port
                           , B2 => n7, ZN => n95);
   U12 : AOI22_X1 port map( A1 => DATA_IN(9), A2 => n4, B1 => DATA_OUT_9_port, 
                           B2 => n7, ZN => n96);
   U11 : AOI22_X1 port map( A1 => DATA_IN(8), A2 => n4, B1 => DATA_OUT_8_port, 
                           B2 => n7, ZN => n97);
   U5 : BUF_X1 port map( A => n1, Z => n7);
   U35 : BUF_X1 port map( A => n1, Z => n6);
   U36 : BUF_X1 port map( A => n1, Z => n8);
   U37 : BUF_X1 port map( A => n2, Z => n4);
   U38 : BUF_X1 port map( A => n2, Z => n3);
   U39 : BUF_X1 port map( A => n2, Z => n5);
   U40 : AND2_X1 port map( A1 => RST, A2 => n9, ZN => n1);
   U41 : AND2_X1 port map( A1 => EN, A2 => RST, ZN => n2);
   U42 : INV_X1 port map( A => EN, ZN => n9);
   U43 : INV_X1 port map( A => n104, ZN => n73);
   U44 : INV_X1 port map( A => n103, ZN => n72);
   U45 : AOI22_X1 port map( A1 => DATA_OUT_2_port, A2 => n8, B1 => DATA_IN(2), 
                           B2 => n5, ZN => n10);
   U46 : INV_X1 port map( A => n10, ZN => n71);
   U47 : INV_X1 port map( A => n102, ZN => n70);
   U48 : INV_X1 port map( A => n101, ZN => n69);
   U49 : INV_X1 port map( A => n100, ZN => n68);
   U50 : INV_X1 port map( A => n99, ZN => n38);
   U51 : INV_X1 port map( A => n98, ZN => n36);
   U52 : INV_X1 port map( A => n97, ZN => n35);
   U53 : INV_X1 port map( A => n96, ZN => n33);
   U54 : INV_X1 port map( A => n95, ZN => n32);
   U55 : INV_X1 port map( A => n94, ZN => n31);
   U56 : INV_X1 port map( A => n93, ZN => n30);
   U57 : INV_X1 port map( A => n92, ZN => n29);
   U58 : INV_X1 port map( A => n91, ZN => n28);
   U59 : INV_X1 port map( A => n90, ZN => n27);
   U60 : INV_X1 port map( A => n89, ZN => n26);
   U61 : INV_X1 port map( A => n88, ZN => n25);
   U62 : INV_X1 port map( A => n87, ZN => n24);
   U63 : INV_X1 port map( A => n86, ZN => n23);
   U64 : INV_X1 port map( A => n85, ZN => n22);
   U65 : INV_X1 port map( A => n84, ZN => n21);
   U66 : INV_X1 port map( A => n83, ZN => n20);
   U67 : INV_X1 port map( A => n82, ZN => n19);
   U68 : INV_X1 port map( A => n81, ZN => n18);
   U69 : INV_X1 port map( A => n80, ZN => n17);
   U70 : INV_X1 port map( A => n79, ZN => n16);
   U71 : INV_X1 port map( A => n78, ZN => n15);
   U72 : INV_X1 port map( A => n77, ZN => n14);
   U73 : INV_X1 port map( A => n76, ZN => n13);
   U74 : INV_X1 port map( A => n75, ZN => n12);
   U75 : INV_X1 port map( A => n74, ZN => n11);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_8 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_8;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, 
      n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, 
      n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, 
      n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377 : 
      std_logic;

begin
   DATA_OUT <= ( DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port );
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n44, CK => CLK, Q => 
                           DATA_OUT_31_port, QN => n_2346);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n45, CK => CLK, Q => 
                           DATA_OUT_30_port, QN => n_2347);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n46, CK => CLK, Q => 
                           DATA_OUT_29_port, QN => n_2348);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n47, CK => CLK, Q => 
                           DATA_OUT_28_port, QN => n_2349);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n48, CK => CLK, Q => 
                           DATA_OUT_27_port, QN => n_2350);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n49, CK => CLK, Q => 
                           DATA_OUT_26_port, QN => n_2351);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n50, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_2352);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n51, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n_2353);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n52, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_2354);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n53, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n_2355);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n54, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n_2356);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n55, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_2357);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n56, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_2358);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n57, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_2359);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n58, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_2360);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n59, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n_2361);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n60, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n_2362);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n61, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n_2363);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n62, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n_2364);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n63, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n_2365);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n64, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n_2366);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n65, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n_2367);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n66, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n_2368);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n67, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n_2369);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n_2370);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n_2371);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT_5_port, QN => n_2372);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_2373);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_2374);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_2375);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_2376);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_2377);
   U3 : BUF_X2 port map( A => n42, Z => n7);
   U4 : BUF_X2 port map( A => n42, Z => n8);
   U5 : BUF_X1 port map( A => n1, Z => n4);
   U6 : BUF_X1 port map( A => n1, Z => n5);
   U7 : BUF_X1 port map( A => n42, Z => n9);
   U8 : BUF_X1 port map( A => n1, Z => n6);
   U9 : AND2_X1 port map( A1 => n2, A2 => n10, ZN => n1);
   U10 : INV_X1 port map( A => n3, ZN => n2);
   U11 : INV_X1 port map( A => RST, ZN => n3);
   U12 : OR2_X1 port map( A1 => EN, A2 => n3, ZN => n10);
   U13 : INV_X1 port map( A => n10, ZN => n42);
   U14 : AOI22_X1 port map( A1 => DATA_OUT_0_port, A2 => n7, B1 => DATA_IN(0), 
                           B2 => n4, ZN => n11);
   U15 : INV_X1 port map( A => n11, ZN => n75);
   U16 : AOI22_X1 port map( A1 => DATA_OUT_1_port, A2 => n7, B1 => DATA_IN(1), 
                           B2 => n4, ZN => n12);
   U17 : INV_X1 port map( A => n12, ZN => n74);
   U18 : AOI22_X1 port map( A1 => DATA_OUT_2_port, A2 => n7, B1 => DATA_IN(2), 
                           B2 => n4, ZN => n13);
   U19 : INV_X1 port map( A => n13, ZN => n73);
   U20 : AOI22_X1 port map( A1 => DATA_OUT_3_port, A2 => n7, B1 => DATA_IN(3), 
                           B2 => n4, ZN => n14);
   U21 : INV_X1 port map( A => n14, ZN => n72);
   U22 : AOI22_X1 port map( A1 => DATA_OUT_4_port, A2 => n7, B1 => DATA_IN(4), 
                           B2 => n4, ZN => n15);
   U23 : INV_X1 port map( A => n15, ZN => n71);
   U24 : AOI22_X1 port map( A1 => DATA_OUT_5_port, A2 => n7, B1 => DATA_IN(5), 
                           B2 => n4, ZN => n16);
   U25 : INV_X1 port map( A => n16, ZN => n70);
   U26 : AOI22_X1 port map( A1 => DATA_OUT_6_port, A2 => n7, B1 => DATA_IN(6), 
                           B2 => n4, ZN => n17);
   U27 : INV_X1 port map( A => n17, ZN => n69);
   U28 : AOI22_X1 port map( A1 => DATA_OUT_7_port, A2 => n7, B1 => DATA_IN(7), 
                           B2 => n4, ZN => n18);
   U29 : INV_X1 port map( A => n18, ZN => n68);
   U30 : AOI22_X1 port map( A1 => DATA_OUT_8_port, A2 => n7, B1 => DATA_IN(8), 
                           B2 => n4, ZN => n19);
   U31 : INV_X1 port map( A => n19, ZN => n67);
   U32 : AOI22_X1 port map( A1 => DATA_OUT_9_port, A2 => n7, B1 => DATA_IN(9), 
                           B2 => n4, ZN => n20);
   U33 : INV_X1 port map( A => n20, ZN => n66);
   U34 : AOI22_X1 port map( A1 => DATA_OUT_10_port, A2 => n7, B1 => DATA_IN(10)
                           , B2 => n4, ZN => n21);
   U35 : INV_X1 port map( A => n21, ZN => n65);
   U36 : AOI22_X1 port map( A1 => DATA_OUT_11_port, A2 => n7, B1 => DATA_IN(11)
                           , B2 => n4, ZN => n22);
   U37 : INV_X1 port map( A => n22, ZN => n64);
   U38 : AOI22_X1 port map( A1 => DATA_OUT_12_port, A2 => n8, B1 => DATA_IN(12)
                           , B2 => n5, ZN => n23);
   U39 : INV_X1 port map( A => n23, ZN => n63);
   U40 : AOI22_X1 port map( A1 => DATA_OUT_13_port, A2 => n8, B1 => DATA_IN(13)
                           , B2 => n5, ZN => n24);
   U41 : INV_X1 port map( A => n24, ZN => n62);
   U42 : AOI22_X1 port map( A1 => DATA_OUT_14_port, A2 => n8, B1 => DATA_IN(14)
                           , B2 => n5, ZN => n25);
   U43 : INV_X1 port map( A => n25, ZN => n61);
   U44 : AOI22_X1 port map( A1 => DATA_OUT_15_port, A2 => n8, B1 => DATA_IN(15)
                           , B2 => n5, ZN => n26);
   U45 : INV_X1 port map( A => n26, ZN => n60);
   U46 : AOI22_X1 port map( A1 => DATA_OUT_16_port, A2 => n8, B1 => DATA_IN(16)
                           , B2 => n5, ZN => n27);
   U47 : INV_X1 port map( A => n27, ZN => n59);
   U48 : AOI22_X1 port map( A1 => DATA_OUT_17_port, A2 => n8, B1 => DATA_IN(17)
                           , B2 => n5, ZN => n28);
   U49 : INV_X1 port map( A => n28, ZN => n58);
   U50 : AOI22_X1 port map( A1 => DATA_OUT_18_port, A2 => n8, B1 => DATA_IN(18)
                           , B2 => n5, ZN => n29);
   U51 : INV_X1 port map( A => n29, ZN => n57);
   U52 : AOI22_X1 port map( A1 => DATA_OUT_19_port, A2 => n8, B1 => DATA_IN(19)
                           , B2 => n5, ZN => n30);
   U53 : INV_X1 port map( A => n30, ZN => n56);
   U54 : AOI22_X1 port map( A1 => DATA_OUT_20_port, A2 => n8, B1 => DATA_IN(20)
                           , B2 => n5, ZN => n31);
   U55 : INV_X1 port map( A => n31, ZN => n55);
   U56 : AOI22_X1 port map( A1 => DATA_OUT_21_port, A2 => n8, B1 => DATA_IN(21)
                           , B2 => n5, ZN => n32);
   U57 : INV_X1 port map( A => n32, ZN => n54);
   U58 : AOI22_X1 port map( A1 => DATA_OUT_22_port, A2 => n8, B1 => DATA_IN(22)
                           , B2 => n5, ZN => n33);
   U59 : INV_X1 port map( A => n33, ZN => n53);
   U60 : AOI22_X1 port map( A1 => DATA_OUT_23_port, A2 => n8, B1 => DATA_IN(23)
                           , B2 => n5, ZN => n34);
   U61 : INV_X1 port map( A => n34, ZN => n52);
   U62 : AOI22_X1 port map( A1 => DATA_OUT_24_port, A2 => n9, B1 => DATA_IN(24)
                           , B2 => n6, ZN => n35);
   U63 : INV_X1 port map( A => n35, ZN => n51);
   U64 : AOI22_X1 port map( A1 => DATA_OUT_25_port, A2 => n9, B1 => DATA_IN(25)
                           , B2 => n6, ZN => n36);
   U65 : INV_X1 port map( A => n36, ZN => n50);
   U66 : AOI22_X1 port map( A1 => DATA_OUT_26_port, A2 => n9, B1 => DATA_IN(26)
                           , B2 => n6, ZN => n37);
   U67 : INV_X1 port map( A => n37, ZN => n49);
   U68 : AOI22_X1 port map( A1 => DATA_OUT_27_port, A2 => n9, B1 => DATA_IN(27)
                           , B2 => n6, ZN => n38);
   U69 : INV_X1 port map( A => n38, ZN => n48);
   U70 : AOI22_X1 port map( A1 => DATA_OUT_28_port, A2 => n9, B1 => DATA_IN(28)
                           , B2 => n6, ZN => n39);
   U71 : INV_X1 port map( A => n39, ZN => n47);
   U72 : AOI22_X1 port map( A1 => DATA_OUT_29_port, A2 => n9, B1 => DATA_IN(29)
                           , B2 => n6, ZN => n40);
   U73 : INV_X1 port map( A => n40, ZN => n46);
   U74 : AOI22_X1 port map( A1 => DATA_OUT_30_port, A2 => n9, B1 => DATA_IN(30)
                           , B2 => n6, ZN => n41);
   U75 : INV_X1 port map( A => n41, ZN => n45);
   U76 : AOI22_X1 port map( A1 => DATA_OUT_31_port, A2 => n9, B1 => DATA_IN(31)
                           , B2 => n6, ZN => n43);
   U77 : INV_X1 port map( A => n43, ZN => n44);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity dlx_cu is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
         EQ_COND, IS_JUMP : out std_logic;  ALU_OPCODE : out std_logic_vector 
         (0 to 3);  DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, IS_JAL, 
         WB_MUX_SEL, RF_WE : out std_logic);

end dlx_cu;

architecture SYN_dlx_cu_hw of dlx_cu is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal aluOpcode1_3_port, aluOpcode1_2_port, aluOpcode1_1_port, 
      aluOpcode1_0_port, aluOpcode_i_3_port, aluOpcode_i_2_port, 
      aluOpcode_i_1_port, aluOpcode_i_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n_2378, 
      n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385 : std_logic;

begin
   
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_3_port, QN => n_2378);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_2_port, QN => n_2379);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_1_port, QN => n_2380);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_0_port, QN => n_2381);
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => aluOpcode1_3_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(0), QN => n_2382);
   aluOpcode2_reg_2_inst : DFFR_X1 port map( D => aluOpcode1_2_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(1), QN => n_2383);
   aluOpcode2_reg_1_inst : DFFR_X1 port map( D => aluOpcode1_1_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(2), QN => n_2384);
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => aluOpcode1_0_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(3), QN => n_2385);
   RF_WE <= '0';
   WB_MUX_SEL <= '0';
   IS_JAL <= '0';
   PC_LATCH_EN <= '0';
   JUMP_EN <= '0';
   LMD_LATCH_EN <= '0';
   DRAM_WE <= '0';
   IS_JUMP <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   SIGNED_IMM <= '0';
   NPC_LATCH_EN <= '0';
   IR_LATCH_EN <= '0';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   U21 : NOR2_X1 port map( A1 => n9, A2 => n8, ZN => n11);
   U22 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => n8);
   U23 : INV_X1 port map( A => IR_IN(10), ZN => n7);
   U24 : AND3_X1 port map( A1 => n44, A2 => n29, A3 => n13, ZN => n1);
   U25 : AND3_X1 port map( A1 => IR_IN(26), A2 => n44, A3 => n29, ZN => n2);
   U26 : NOR2_X1 port map( A1 => IR_IN(7), A2 => IR_IN(4), ZN => n5);
   U27 : INV_X1 port map( A => IR_IN(9), ZN => n6);
   U28 : INV_X1 port map( A => IR_IN(8), ZN => n3);
   U29 : INV_X1 port map( A => IR_IN(6), ZN => n4);
   U30 : NAND3_X1 port map( A1 => n5, A2 => n4, A3 => n3, ZN => n9);
   U31 : NAND2_X1 port map( A1 => IR_IN(5), A2 => n11, ZN => n48);
   U32 : NOR2_X1 port map( A1 => IR_IN(3), A2 => n48, ZN => n12);
   U33 : INV_X1 port map( A => IR_IN(2), ZN => n59);
   U34 : NAND2_X1 port map( A1 => IR_IN(1), A2 => n59, ZN => n35);
   U35 : INV_X1 port map( A => IR_IN(3), ZN => n50);
   U36 : INV_X1 port map( A => IR_IN(5), ZN => n10);
   U37 : NAND4_X1 port map( A1 => IR_IN(2), A2 => n11, A3 => n50, A4 => n10, ZN
                           => n39);
   U38 : INV_X1 port map( A => n39, ZN => n61);
   U39 : AOI22_X1 port map( A1 => n12, A2 => n35, B1 => IR_IN(1), B2 => n61, ZN
                           => n26);
   U40 : INV_X1 port map( A => IR_IN(27), ZN => n44);
   U41 : INV_X1 port map( A => IR_IN(31), ZN => n29);
   U42 : INV_X1 port map( A => IR_IN(30), ZN => n23);
   U43 : INV_X1 port map( A => IR_IN(29), ZN => n56);
   U44 : NAND2_X1 port map( A1 => n23, A2 => n56, ZN => n31);
   U45 : NOR3_X1 port map( A1 => IR_IN(26), A2 => IR_IN(28), A3 => n31, ZN => 
                           n13);
   U46 : INV_X1 port map( A => IR_IN(0), ZN => n49);
   U47 : NAND2_X1 port map( A1 => n1, A2 => n49, ZN => n34);
   U48 : INV_X1 port map( A => IR_IN(28), ZN => n16);
   U49 : NAND3_X1 port map( A1 => IR_IN(29), A2 => IR_IN(30), A3 => n2, ZN => 
                           n65);
   U50 : INV_X1 port map( A => IR_IN(1), ZN => n36);
   U51 : NOR3_X1 port map( A1 => n48, A2 => n50, A3 => n49, ZN => n14);
   U52 : NAND3_X1 port map( A1 => n1, A2 => n36, A3 => n14, ZN => n58);
   U53 : OAI22_X1 port map( A1 => n16, A2 => n65, B1 => n59, B2 => n58, ZN => 
                           n15);
   U54 : INV_X1 port map( A => n15, ZN => n55);
   U55 : INV_X1 port map( A => IR_IN(26), ZN => n30);
   U56 : NAND3_X1 port map( A1 => IR_IN(28), A2 => n30, A3 => n29, ZN => n32);
   U57 : MUX2_X1 port map( A => IR_IN(28), B => n30, S => IR_IN(29), Z => n17);
   U58 : NAND2_X1 port map( A1 => IR_IN(27), A2 => n16, ZN => n27);
   U59 : INV_X1 port map( A => n27, ZN => n18);
   U60 : AOI22_X1 port map( A1 => n17, A2 => n44, B1 => n18, B2 => n56, ZN => 
                           n20);
   U61 : NAND2_X1 port map( A1 => n18, A2 => IR_IN(26), ZN => n19);
   U62 : MUX2_X1 port map( A => n20, B => n19, S => IR_IN(31), Z => n21);
   U63 : OAI21_X1 port map( B1 => n32, B2 => n56, A => n21, ZN => n24);
   U64 : INV_X1 port map( A => n32, ZN => n45);
   U65 : NAND3_X1 port map( A1 => IR_IN(30), A2 => n45, A3 => n56, ZN => n64);
   U66 : INV_X1 port map( A => n64, ZN => n22);
   U67 : AOI22_X1 port map( A1 => n24, A2 => n23, B1 => n22, B2 => IR_IN(27), 
                           ZN => n25);
   U68 : OAI211_X1 port map( C1 => n26, C2 => n34, A => n55, B => n25, ZN => 
                           aluOpcode_i_0_port);
   U69 : NOR3_X1 port map( A1 => IR_IN(30), A2 => n56, A3 => n27, ZN => n28);
   U70 : NAND3_X1 port map( A1 => n30, A2 => n29, A3 => n28, ZN => n43);
   U71 : INV_X1 port map( A => n31, ZN => n33);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n32, ZN => n41);
   U73 : INV_X1 port map( A => n34, ZN => n62);
   U74 : INV_X1 port map( A => n35, ZN => n37);
   U75 : AOI22_X1 port map( A1 => n37, A2 => n50, B1 => IR_IN(2), B2 => n36, ZN
                           => n38);
   U76 : OAI22_X1 port map( A1 => IR_IN(1), A2 => n39, B1 => n38, B2 => n48, ZN
                           => n40);
   U77 : AOI22_X1 port map( A1 => n41, A2 => n44, B1 => n62, B2 => n40, ZN => 
                           n42);
   U78 : NAND3_X1 port map( A1 => n55, A2 => n43, A3 => n42, ZN => 
                           aluOpcode_i_1_port);
   U79 : AOI22_X1 port map( A1 => n2, A2 => IR_IN(28), B1 => IR_IN(27), B2 => 
                           n45, ZN => n47);
   U80 : NAND2_X1 port map( A1 => n45, A2 => n44, ZN => n46);
   U81 : MUX2_X1 port map( A => n47, B => n46, S => IR_IN(30), Z => n57);
   U82 : INV_X1 port map( A => n48, ZN => n53);
   U83 : NAND2_X1 port map( A1 => n50, A2 => n49, ZN => n51);
   U84 : XOR2_X1 port map( A => n51, B => IR_IN(1), Z => n52);
   U85 : NAND4_X1 port map( A1 => n53, A2 => IR_IN(2), A3 => n1, A4 => n52, ZN 
                           => n54);
   U86 : OAI211_X1 port map( C1 => n57, C2 => n56, A => n55, B => n54, ZN => 
                           aluOpcode_i_2_port);
   U87 : INV_X1 port map( A => n58, ZN => n60);
   U88 : AOI22_X1 port map( A1 => n62, A2 => n61, B1 => n60, B2 => n59, ZN => 
                           n63);
   U89 : OAI211_X1 port map( C1 => IR_IN(28), C2 => n65, A => n64, B => n63, ZN
                           => aluOpcode_i_3_port);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 is

   port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
         EQ_COND, IS_JUMP : in std_logic;  ALU_OPCODE : in std_logic_vector (0 
         to 3);  JUMP_EN, PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE : in std_logic
         ;  D_ADDR : out std_logic_vector (5 downto 0);  D_DATA_IN : out 
         std_logic_vector (31 downto 0);  D_DATA_OUT, PC_IN : in 
         std_logic_vector (31 downto 0);  PC_BUS : out std_logic_vector (31 
         downto 0));

end DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64;

architecture SYN_STRUCTURE of 
   DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 is

   component ALU_N32
      port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26
      port( NOT_EXT_IMM : in std_logic_vector (25 downto 0);  SIGNED_IMM, 
            IS_JUMP : in std_logic;  EXT_IMM : out std_logic_vector (31 downto 
            0));
   end component;
   
   component REGISTER_FILE_NBIT32_NREG32
      port( CLK, RST, EN, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component ADDER_N32
      port( CURR_ADDR : in std_logic_vector (31 downto 0);  NEXT_ADDR : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT5_1
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT5_0
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component MUX21
      port( A, B, SEL : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component BRANCHING_UNIT_N32
      port( CLK, RST : in std_logic;  Reg_A : in std_logic_vector (31 downto 0)
            ;  EQ_cond, IS_JUMP : in std_logic;  branch_taken : out std_logic);
   end component;
   
   component REG_GENERIC_NBIT32_1
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_2
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_3
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT5_1
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 
            downto 0);  DATA_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component REG_GENERIC_NBIT5_2
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 
            downto 0);  DATA_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component REG_GENERIC_NBIT5_0
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 
            downto 0);  DATA_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component REG_GENERIC_NBIT26
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (25 
            downto 0);  DATA_OUT : out std_logic_vector (25 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_4
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_5
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_6
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_7
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_8
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, D_ADDR_5_port, D_ADDR_4_port, 
      D_ADDR_3_port, D_ADDR_2_port, D_ADDR_1_port, D_ADDR_0_port, 
      PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, current_PC_31_port, 
      current_PC_30_port, current_PC_29_port, current_PC_28_port, 
      current_PC_27_port, current_PC_26_port, current_PC_25_port, 
      current_PC_24_port, current_PC_23_port, current_PC_22_port, 
      current_PC_21_port, current_PC_20_port, current_PC_19_port, 
      current_PC_18_port, current_PC_17_port, current_PC_16_port, 
      current_PC_15_port, current_PC_14_port, current_PC_13_port, 
      current_PC_12_port, current_PC_11_port, current_PC_10_port, 
      current_PC_9_port, current_PC_8_port, current_PC_7_port, 
      current_PC_6_port, current_PC_5_port, current_PC_4_port, 
      current_PC_3_port, current_PC_2_port, current_PC_1_port, 
      current_PC_0_port, current_PC1_31_port, current_PC1_30_port, 
      current_PC1_29_port, current_PC1_28_port, current_PC1_27_port, 
      current_PC1_26_port, current_PC1_25_port, current_PC1_24_port, 
      current_PC1_23_port, current_PC1_22_port, current_PC1_21_port, 
      current_PC1_20_port, current_PC1_19_port, current_PC1_18_port, 
      current_PC1_17_port, current_PC1_16_port, current_PC1_15_port, 
      current_PC1_14_port, current_PC1_13_port, current_PC1_12_port, 
      current_PC1_11_port, current_PC1_10_port, current_PC1_9_port, 
      current_PC1_8_port, current_PC1_7_port, current_PC1_6_port, 
      current_PC1_5_port, current_PC1_4_port, current_PC1_3_port, 
      current_PC1_2_port, current_PC1_1_port, current_PC1_0_port, 
      current_PC2_31_port, current_PC2_30_port, current_PC2_29_port, 
      current_PC2_28_port, current_PC2_27_port, current_PC2_26_port, 
      current_PC2_25_port, current_PC2_24_port, current_PC2_23_port, 
      current_PC2_22_port, current_PC2_21_port, current_PC2_20_port, 
      current_PC2_19_port, current_PC2_18_port, current_PC2_17_port, 
      current_PC2_16_port, current_PC2_15_port, current_PC2_14_port, 
      current_PC2_13_port, current_PC2_12_port, current_PC2_11_port, 
      current_PC2_10_port, current_PC2_9_port, current_PC2_8_port, 
      current_PC2_7_port, current_PC2_6_port, current_PC2_5_port, 
      current_PC2_4_port, current_PC2_3_port, current_PC2_2_port, 
      current_PC2_1_port, current_PC2_0_port, current_PC3_31_port, 
      current_PC3_30_port, current_PC3_29_port, current_PC3_28_port, 
      current_PC3_27_port, current_PC3_26_port, current_PC3_25_port, 
      current_PC3_24_port, current_PC3_23_port, current_PC3_22_port, 
      current_PC3_21_port, current_PC3_20_port, current_PC3_19_port, 
      current_PC3_18_port, current_PC3_17_port, current_PC3_16_port, 
      current_PC3_15_port, current_PC3_14_port, current_PC3_13_port, 
      current_PC3_12_port, current_PC3_11_port, current_PC3_10_port, 
      current_PC3_9_port, current_PC3_8_port, current_PC3_7_port, 
      current_PC3_6_port, current_PC3_5_port, current_PC3_4_port, 
      current_PC3_3_port, current_PC3_2_port, current_PC3_1_port, 
      current_PC3_0_port, next_NPC_31_port, next_NPC_30_port, next_NPC_29_port,
      next_NPC_28_port, next_NPC_27_port, next_NPC_26_port, next_NPC_25_port, 
      next_NPC_24_port, next_NPC_23_port, next_NPC_22_port, next_NPC_21_port, 
      next_NPC_20_port, next_NPC_19_port, next_NPC_18_port, next_NPC_17_port, 
      next_NPC_16_port, next_NPC_15_port, next_NPC_14_port, next_NPC_13_port, 
      next_NPC_12_port, next_NPC_11_port, next_NPC_10_port, next_NPC_9_port, 
      next_NPC_8_port, next_NPC_7_port, next_NPC_6_port, next_NPC_5_port, 
      next_NPC_4_port, next_NPC_3_port, next_NPC_2_port, next_NPC_1_port, 
      next_NPC_0_port, current_NPC_31_port, current_NPC_30_port, 
      current_NPC_29_port, current_NPC_28_port, current_NPC_27_port, 
      current_NPC_26_port, current_NPC_25_port, current_NPC_24_port, 
      current_NPC_23_port, current_NPC_22_port, current_NPC_21_port, 
      current_NPC_20_port, current_NPC_19_port, current_NPC_18_port, 
      current_NPC_17_port, current_NPC_16_port, current_NPC_15_port, 
      current_NPC_14_port, current_NPC_13_port, current_NPC_12_port, 
      current_NPC_11_port, current_NPC_10_port, current_NPC_9_port, 
      current_NPC_8_port, current_NPC_7_port, current_NPC_6_port, 
      current_NPC_5_port, current_NPC_4_port, current_NPC_3_port, 
      current_NPC_2_port, current_NPC_1_port, current_NPC_0_port, 
      current_IW_25_port, current_IW_24_port, current_IW_23_port, 
      current_IW_22_port, current_IW_21_port, current_IW_20_port, 
      current_IW_19_port, current_IW_18_port, current_IW_17_port, 
      current_IW_16_port, current_IW_15_port, current_IW_14_port, 
      current_IW_13_port, current_IW_12_port, current_IW_11_port, 
      current_IW_10_port, current_IW_9_port, current_IW_8_port, 
      current_IW_7_port, current_IW_6_port, current_IW_5_port, 
      current_IW_4_port, current_IW_3_port, current_IW_2_port, 
      current_IW_1_port, current_IW_0_port, IMM_IN_25_port, IMM_IN_24_port, 
      IMM_IN_23_port, IMM_IN_22_port, IMM_IN_21_port, IMM_IN_20_port, 
      IMM_IN_19_port, IMM_IN_18_port, IMM_IN_17_port, IMM_IN_16_port, 
      IMM_IN_15_port, IMM_IN_14_port, IMM_IN_13_port, IMM_IN_12_port, 
      IMM_IN_11_port, IMM_IN_10_port, IMM_IN_9_port, IMM_IN_8_port, 
      IMM_IN_7_port, IMM_IN_6_port, IMM_IN_5_port, IMM_IN_4_port, IMM_IN_3_port
      , IMM_IN_2_port, IMM_IN_1_port, IMM_IN_0_port, WB1_IN_4_port, 
      WB1_IN_3_port, WB1_IN_2_port, WB1_IN_1_port, WB1_IN_0_port, WB2_IN_4_port
      , WB2_IN_3_port, WB2_IN_2_port, WB2_IN_1_port, WB2_IN_0_port, 
      WB2_OUT_4_port, WB2_OUT_3_port, WB2_OUT_2_port, WB2_OUT_1_port, 
      WB2_OUT_0_port, WB3_OUT_4_port, WB3_OUT_3_port, WB3_OUT_2_port, 
      WB3_OUT_1_port, WB3_OUT_0_port, next_ALU_OUT_31_port, 
      next_ALU_OUT_30_port, next_ALU_OUT_29_port, next_ALU_OUT_28_port, 
      next_ALU_OUT_27_port, next_ALU_OUT_26_port, next_ALU_OUT_25_port, 
      next_ALU_OUT_24_port, next_ALU_OUT_23_port, next_ALU_OUT_22_port, 
      next_ALU_OUT_21_port, next_ALU_OUT_20_port, next_ALU_OUT_19_port, 
      next_ALU_OUT_18_port, next_ALU_OUT_17_port, next_ALU_OUT_16_port, 
      next_ALU_OUT_15_port, next_ALU_OUT_14_port, next_ALU_OUT_13_port, 
      next_ALU_OUT_12_port, next_ALU_OUT_11_port, next_ALU_OUT_10_port, 
      next_ALU_OUT_9_port, next_ALU_OUT_8_port, next_ALU_OUT_7_port, 
      next_ALU_OUT_6_port, next_ALU_OUT_5_port, next_ALU_OUT_4_port, 
      next_ALU_OUT_3_port, next_ALU_OUT_2_port, next_ALU_OUT_1_port, 
      next_ALU_OUT_0_port, current_ALU_OUT_31_port, current_ALU_OUT_30_port, 
      current_ALU_OUT_29_port, current_ALU_OUT_28_port, current_ALU_OUT_27_port
      , current_ALU_OUT_26_port, current_ALU_OUT_25_port, 
      current_ALU_OUT_24_port, current_ALU_OUT_23_port, current_ALU_OUT_22_port
      , current_ALU_OUT_21_port, current_ALU_OUT_20_port, 
      current_ALU_OUT_19_port, current_ALU_OUT_18_port, current_ALU_OUT_17_port
      , current_ALU_OUT_16_port, current_ALU_OUT_15_port, 
      current_ALU_OUT_14_port, current_ALU_OUT_13_port, current_ALU_OUT_12_port
      , current_ALU_OUT_11_port, current_ALU_OUT_10_port, 
      current_ALU_OUT_9_port, current_ALU_OUT_8_port, current_ALU_OUT_7_port, 
      current_ALU_OUT_6_port, B_OUT_31_port, B_OUT_30_port, B_OUT_29_port, 
      B_OUT_28_port, B_OUT_27_port, B_OUT_26_port, B_OUT_25_port, B_OUT_24_port
      , B_OUT_23_port, B_OUT_22_port, B_OUT_21_port, B_OUT_20_port, 
      B_OUT_19_port, B_OUT_18_port, B_OUT_17_port, B_OUT_16_port, B_OUT_15_port
      , B_OUT_14_port, B_OUT_13_port, B_OUT_12_port, B_OUT_11_port, 
      B_OUT_10_port, B_OUT_9_port, B_OUT_8_port, B_OUT_7_port, B_OUT_6_port, 
      B_OUT_5_port, B_OUT_4_port, B_OUT_3_port, B_OUT_2_port, B_OUT_1_port, 
      B_OUT_0_port, current_ALU_OUT2_31_port, current_ALU_OUT2_30_port, 
      current_ALU_OUT2_29_port, current_ALU_OUT2_28_port, 
      current_ALU_OUT2_27_port, current_ALU_OUT2_26_port, 
      current_ALU_OUT2_25_port, current_ALU_OUT2_24_port, 
      current_ALU_OUT2_23_port, current_ALU_OUT2_22_port, 
      current_ALU_OUT2_21_port, current_ALU_OUT2_20_port, 
      current_ALU_OUT2_19_port, current_ALU_OUT2_18_port, 
      current_ALU_OUT2_17_port, current_ALU_OUT2_16_port, 
      current_ALU_OUT2_15_port, current_ALU_OUT2_14_port, 
      current_ALU_OUT2_13_port, current_ALU_OUT2_12_port, 
      current_ALU_OUT2_11_port, current_ALU_OUT2_10_port, 
      current_ALU_OUT2_9_port, current_ALU_OUT2_8_port, current_ALU_OUT2_7_port
      , current_ALU_OUT2_6_port, current_ALU_OUT2_5_port, 
      current_ALU_OUT2_4_port, current_ALU_OUT2_3_port, current_ALU_OUT2_2_port
      , current_ALU_OUT2_1_port, current_ALU_OUT2_0_port, A_OUT_31_port, 
      A_OUT_30_port, A_OUT_29_port, A_OUT_28_port, A_OUT_27_port, A_OUT_26_port
      , A_OUT_25_port, A_OUT_24_port, A_OUT_23_port, A_OUT_22_port, 
      A_OUT_21_port, A_OUT_20_port, A_OUT_19_port, A_OUT_18_port, A_OUT_17_port
      , A_OUT_16_port, A_OUT_15_port, A_OUT_14_port, A_OUT_13_port, 
      A_OUT_12_port, A_OUT_11_port, A_OUT_10_port, A_OUT_9_port, A_OUT_8_port, 
      A_OUT_7_port, A_OUT_6_port, A_OUT_5_port, A_OUT_4_port, A_OUT_3_port, 
      A_OUT_2_port, A_OUT_1_port, A_OUT_0_port, branch_taken, PC_MUX_SEL, 
      ALU_OP1_31_port, ALU_OP1_30_port, ALU_OP1_29_port, ALU_OP1_28_port, 
      ALU_OP1_27_port, ALU_OP1_26_port, ALU_OP1_25_port, ALU_OP1_24_port, 
      ALU_OP1_23_port, ALU_OP1_22_port, ALU_OP1_21_port, ALU_OP1_20_port, 
      ALU_OP1_19_port, ALU_OP1_18_port, ALU_OP1_17_port, ALU_OP1_16_port, 
      ALU_OP1_15_port, ALU_OP1_14_port, ALU_OP1_13_port, ALU_OP1_12_port, 
      ALU_OP1_11_port, ALU_OP1_10_port, ALU_OP1_9_port, ALU_OP1_8_port, 
      ALU_OP1_7_port, ALU_OP1_6_port, ALU_OP1_5_port, ALU_OP1_4_port, 
      ALU_OP1_3_port, ALU_OP1_2_port, ALU_OP1_1_port, ALU_OP1_0_port, 
      IMM_OUT_31_port, IMM_OUT_30_port, IMM_OUT_29_port, IMM_OUT_28_port, 
      IMM_OUT_27_port, IMM_OUT_26_port, IMM_OUT_25_port, IMM_OUT_24_port, 
      IMM_OUT_23_port, IMM_OUT_22_port, IMM_OUT_21_port, IMM_OUT_20_port, 
      IMM_OUT_19_port, IMM_OUT_18_port, IMM_OUT_17_port, IMM_OUT_16_port, 
      IMM_OUT_15_port, IMM_OUT_14_port, IMM_OUT_13_port, IMM_OUT_12_port, 
      IMM_OUT_11_port, IMM_OUT_10_port, IMM_OUT_9_port, IMM_OUT_8_port, 
      IMM_OUT_7_port, IMM_OUT_6_port, IMM_OUT_5_port, IMM_OUT_4_port, 
      IMM_OUT_3_port, IMM_OUT_2_port, IMM_OUT_1_port, IMM_OUT_0_port, 
      ALU_OP2_31_port, ALU_OP2_30_port, ALU_OP2_29_port, ALU_OP2_28_port, 
      ALU_OP2_27_port, ALU_OP2_26_port, ALU_OP2_25_port, ALU_OP2_24_port, 
      ALU_OP2_23_port, ALU_OP2_22_port, ALU_OP2_21_port, ALU_OP2_20_port, 
      ALU_OP2_19_port, ALU_OP2_18_port, ALU_OP2_17_port, ALU_OP2_16_port, 
      ALU_OP2_15_port, ALU_OP2_14_port, ALU_OP2_13_port, ALU_OP2_12_port, 
      ALU_OP2_11_port, ALU_OP2_10_port, ALU_OP2_9_port, ALU_OP2_8_port, 
      ALU_OP2_7_port, ALU_OP2_6_port, ALU_OP2_5_port, ALU_OP2_4_port, 
      ALU_OP2_3_port, ALU_OP2_2_port, ALU_OP2_1_port, ALU_OP2_0_port, 
      OUT_MUX_DATA_31_port, OUT_MUX_DATA_30_port, OUT_MUX_DATA_29_port, 
      OUT_MUX_DATA_28_port, OUT_MUX_DATA_27_port, OUT_MUX_DATA_26_port, 
      OUT_MUX_DATA_25_port, OUT_MUX_DATA_24_port, OUT_MUX_DATA_23_port, 
      OUT_MUX_DATA_22_port, OUT_MUX_DATA_21_port, OUT_MUX_DATA_20_port, 
      OUT_MUX_DATA_19_port, OUT_MUX_DATA_18_port, OUT_MUX_DATA_17_port, 
      OUT_MUX_DATA_16_port, OUT_MUX_DATA_15_port, OUT_MUX_DATA_14_port, 
      OUT_MUX_DATA_13_port, OUT_MUX_DATA_12_port, OUT_MUX_DATA_11_port, 
      OUT_MUX_DATA_10_port, OUT_MUX_DATA_9_port, OUT_MUX_DATA_8_port, 
      OUT_MUX_DATA_7_port, OUT_MUX_DATA_6_port, OUT_MUX_DATA_5_port, 
      OUT_MUX_DATA_4_port, OUT_MUX_DATA_3_port, OUT_MUX_DATA_2_port, 
      OUT_MUX_DATA_1_port, OUT_MUX_DATA_0_port, WB_DATA_31_port, 
      WB_DATA_30_port, WB_DATA_29_port, WB_DATA_28_port, WB_DATA_27_port, 
      WB_DATA_26_port, WB_DATA_25_port, WB_DATA_24_port, WB_DATA_23_port, 
      WB_DATA_22_port, WB_DATA_21_port, WB_DATA_20_port, WB_DATA_19_port, 
      WB_DATA_18_port, WB_DATA_17_port, WB_DATA_16_port, WB_DATA_15_port, 
      WB_DATA_14_port, WB_DATA_13_port, WB_DATA_12_port, WB_DATA_11_port, 
      WB_DATA_10_port, WB_DATA_9_port, WB_DATA_8_port, WB_DATA_7_port, 
      WB_DATA_6_port, WB_DATA_5_port, WB_DATA_4_port, WB_DATA_3_port, 
      WB_DATA_2_port, WB_DATA_1_port, WB_DATA_0_port, WB_ADDR_4_port, 
      WB_ADDR_3_port, WB_ADDR_2_port, WB_ADDR_1_port, WB_ADDR_0_port, n1, n2, 
      n3, n4, n5, n6, n7, n8, n9, n_2386, n_2387, n_2388, n_2389, n_2390, 
      n_2391 : std_logic;

begin
   D_ADDR <= ( D_ADDR_5_port, D_ADDR_4_port, D_ADDR_3_port, D_ADDR_2_port, 
      D_ADDR_1_port, D_ADDR_0_port );
   PC_BUS <= ( PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U3 : CLKBUF_X1 port map( A => B_OUT_4_port, Z => n1);
   U4 : CLKBUF_X1 port map( A => B_OUT_3_port, Z => n2);
   U5 : AND2_X1 port map( A1 => PC_BUS_0_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_0_port);
   U6 : AND2_X1 port map( A1 => PC_BUS_1_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_1_port);
   U7 : AND2_X1 port map( A1 => PC_BUS_2_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_2_port);
   U8 : AND2_X1 port map( A1 => PC_BUS_3_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_3_port);
   U9 : AND2_X1 port map( A1 => PC_BUS_4_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_4_port);
   U10 : AND2_X1 port map( A1 => PC_BUS_5_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_5_port);
   U11 : AND2_X1 port map( A1 => PC_BUS_6_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_6_port);
   U12 : AND2_X1 port map( A1 => PC_BUS_7_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_7_port);
   U13 : AND2_X1 port map( A1 => PC_BUS_8_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_8_port);
   U14 : AND2_X1 port map( A1 => PC_BUS_10_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_10_port);
   U15 : AND2_X1 port map( A1 => PC_BUS_11_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_11_port);
   U16 : AND2_X1 port map( A1 => PC_BUS_12_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_12_port);
   U17 : AND2_X1 port map( A1 => PC_BUS_13_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_13_port);
   U18 : AND2_X1 port map( A1 => PC_BUS_14_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_14_port);
   U19 : AND2_X1 port map( A1 => PC_BUS_15_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_15_port);
   U20 : AND2_X1 port map( A1 => PC_BUS_16_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_16_port);
   U21 : AND2_X1 port map( A1 => PC_BUS_17_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_17_port);
   U22 : AND2_X1 port map( A1 => PC_BUS_18_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_18_port);
   U23 : AND2_X1 port map( A1 => PC_BUS_19_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_19_port);
   U24 : AND2_X1 port map( A1 => PC_BUS_20_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_20_port);
   U25 : AND2_X1 port map( A1 => PC_BUS_21_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_21_port);
   U26 : AND2_X1 port map( A1 => PC_BUS_22_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_22_port);
   U27 : AND2_X1 port map( A1 => PC_BUS_23_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_23_port);
   U28 : AND2_X1 port map( A1 => PC_BUS_24_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_24_port);
   U29 : AND2_X1 port map( A1 => PC_BUS_25_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_25_port);
   U30 : AND2_X1 port map( A1 => PC_BUS_26_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_26_port);
   U31 : AND2_X1 port map( A1 => PC_BUS_27_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_27_port);
   U32 : AND2_X1 port map( A1 => PC_BUS_28_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_28_port);
   U33 : AND2_X1 port map( A1 => PC_BUS_29_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_29_port);
   U34 : AND2_X1 port map( A1 => PC_BUS_30_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_30_port);
   U35 : AND2_X1 port map( A1 => PC_LATCH_EN, A2 => PC_BUS_9_port, ZN => 
                           current_PC_9_port);
   U36 : AND2_X1 port map( A1 => PC_BUS_31_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_31_port);
   U37 : CLKBUF_X1 port map( A => D_ADDR_0_port, Z => n3);
   U38 : CLKBUF_X1 port map( A => D_ADDR_1_port, Z => n4);
   U39 : CLKBUF_X1 port map( A => D_ADDR_2_port, Z => n5);
   U40 : CLKBUF_X1 port map( A => D_ADDR_3_port, Z => n6);
   U41 : CLKBUF_X1 port map( A => D_ADDR_4_port, Z => n7);
   U42 : CLKBUF_X1 port map( A => D_ADDR_5_port, Z => n8);
   U43 : CLKBUF_X1 port map( A => B_OUT_1_port, Z => n9);
   PC_REG : REG_GENERIC_NBIT32_8 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => PC_IN(31), DATA_IN(30) 
                           => PC_IN(30), DATA_IN(29) => PC_IN(29), DATA_IN(28) 
                           => PC_IN(28), DATA_IN(27) => PC_IN(27), DATA_IN(26) 
                           => PC_IN(26), DATA_IN(25) => PC_IN(25), DATA_IN(24) 
                           => PC_IN(24), DATA_IN(23) => PC_IN(23), DATA_IN(22) 
                           => PC_IN(22), DATA_IN(21) => PC_IN(21), DATA_IN(20) 
                           => PC_IN(20), DATA_IN(19) => PC_IN(19), DATA_IN(18) 
                           => PC_IN(18), DATA_IN(17) => PC_IN(17), DATA_IN(16) 
                           => PC_IN(16), DATA_IN(15) => PC_IN(15), DATA_IN(14) 
                           => PC_IN(14), DATA_IN(13) => PC_IN(13), DATA_IN(12) 
                           => PC_IN(12), DATA_IN(11) => PC_IN(11), DATA_IN(10) 
                           => PC_IN(10), DATA_IN(9) => PC_IN(9), DATA_IN(8) => 
                           PC_IN(8), DATA_IN(7) => PC_IN(7), DATA_IN(6) => 
                           PC_IN(6), DATA_IN(5) => PC_IN(5), DATA_IN(4) => 
                           PC_IN(4), DATA_IN(3) => PC_IN(3), DATA_IN(2) => 
                           PC_IN(2), DATA_IN(1) => PC_IN(1), DATA_IN(0) => 
                           PC_IN(0), DATA_OUT(31) => current_PC1_31_port, 
                           DATA_OUT(30) => current_PC1_30_port, DATA_OUT(29) =>
                           current_PC1_29_port, DATA_OUT(28) => 
                           current_PC1_28_port, DATA_OUT(27) => 
                           current_PC1_27_port, DATA_OUT(26) => 
                           current_PC1_26_port, DATA_OUT(25) => 
                           current_PC1_25_port, DATA_OUT(24) => 
                           current_PC1_24_port, DATA_OUT(23) => 
                           current_PC1_23_port, DATA_OUT(22) => 
                           current_PC1_22_port, DATA_OUT(21) => 
                           current_PC1_21_port, DATA_OUT(20) => 
                           current_PC1_20_port, DATA_OUT(19) => 
                           current_PC1_19_port, DATA_OUT(18) => 
                           current_PC1_18_port, DATA_OUT(17) => 
                           current_PC1_17_port, DATA_OUT(16) => 
                           current_PC1_16_port, DATA_OUT(15) => 
                           current_PC1_15_port, DATA_OUT(14) => 
                           current_PC1_14_port, DATA_OUT(13) => 
                           current_PC1_13_port, DATA_OUT(12) => 
                           current_PC1_12_port, DATA_OUT(11) => 
                           current_PC1_11_port, DATA_OUT(10) => 
                           current_PC1_10_port, DATA_OUT(9) => 
                           current_PC1_9_port, DATA_OUT(8) => 
                           current_PC1_8_port, DATA_OUT(7) => 
                           current_PC1_7_port, DATA_OUT(6) => 
                           current_PC1_6_port, DATA_OUT(5) => 
                           current_PC1_5_port, DATA_OUT(4) => 
                           current_PC1_4_port, DATA_OUT(3) => 
                           current_PC1_3_port, DATA_OUT(2) => 
                           current_PC1_2_port, DATA_OUT(1) => 
                           current_PC1_1_port, DATA_OUT(0) => 
                           current_PC1_0_port);
   PC2_REG : REG_GENERIC_NBIT32_7 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => current_PC1_31_port, 
                           DATA_IN(30) => current_PC1_30_port, DATA_IN(29) => 
                           current_PC1_29_port, DATA_IN(28) => 
                           current_PC1_28_port, DATA_IN(27) => 
                           current_PC1_27_port, DATA_IN(26) => 
                           current_PC1_26_port, DATA_IN(25) => 
                           current_PC1_25_port, DATA_IN(24) => 
                           current_PC1_24_port, DATA_IN(23) => 
                           current_PC1_23_port, DATA_IN(22) => 
                           current_PC1_22_port, DATA_IN(21) => 
                           current_PC1_21_port, DATA_IN(20) => 
                           current_PC1_20_port, DATA_IN(19) => 
                           current_PC1_19_port, DATA_IN(18) => 
                           current_PC1_18_port, DATA_IN(17) => 
                           current_PC1_17_port, DATA_IN(16) => 
                           current_PC1_16_port, DATA_IN(15) => 
                           current_PC1_15_port, DATA_IN(14) => 
                           current_PC1_14_port, DATA_IN(13) => 
                           current_PC1_13_port, DATA_IN(12) => 
                           current_PC1_12_port, DATA_IN(11) => 
                           current_PC1_11_port, DATA_IN(10) => 
                           current_PC1_10_port, DATA_IN(9) => 
                           current_PC1_9_port, DATA_IN(8) => current_PC1_8_port
                           , DATA_IN(7) => current_PC1_7_port, DATA_IN(6) => 
                           current_PC1_6_port, DATA_IN(5) => current_PC1_5_port
                           , DATA_IN(4) => current_PC1_4_port, DATA_IN(3) => 
                           current_PC1_3_port, DATA_IN(2) => current_PC1_2_port
                           , DATA_IN(1) => current_PC1_1_port, DATA_IN(0) => 
                           current_PC1_0_port, DATA_OUT(31) => 
                           current_PC2_31_port, DATA_OUT(30) => 
                           current_PC2_30_port, DATA_OUT(29) => 
                           current_PC2_29_port, DATA_OUT(28) => 
                           current_PC2_28_port, DATA_OUT(27) => 
                           current_PC2_27_port, DATA_OUT(26) => 
                           current_PC2_26_port, DATA_OUT(25) => 
                           current_PC2_25_port, DATA_OUT(24) => 
                           current_PC2_24_port, DATA_OUT(23) => 
                           current_PC2_23_port, DATA_OUT(22) => 
                           current_PC2_22_port, DATA_OUT(21) => 
                           current_PC2_21_port, DATA_OUT(20) => 
                           current_PC2_20_port, DATA_OUT(19) => 
                           current_PC2_19_port, DATA_OUT(18) => 
                           current_PC2_18_port, DATA_OUT(17) => 
                           current_PC2_17_port, DATA_OUT(16) => 
                           current_PC2_16_port, DATA_OUT(15) => 
                           current_PC2_15_port, DATA_OUT(14) => 
                           current_PC2_14_port, DATA_OUT(13) => 
                           current_PC2_13_port, DATA_OUT(12) => 
                           current_PC2_12_port, DATA_OUT(11) => 
                           current_PC2_11_port, DATA_OUT(10) => 
                           current_PC2_10_port, DATA_OUT(9) => 
                           current_PC2_9_port, DATA_OUT(8) => 
                           current_PC2_8_port, DATA_OUT(7) => 
                           current_PC2_7_port, DATA_OUT(6) => 
                           current_PC2_6_port, DATA_OUT(5) => 
                           current_PC2_5_port, DATA_OUT(4) => 
                           current_PC2_4_port, DATA_OUT(3) => 
                           current_PC2_3_port, DATA_OUT(2) => 
                           current_PC2_2_port, DATA_OUT(1) => 
                           current_PC2_1_port, DATA_OUT(0) => 
                           current_PC2_0_port);
   PC3_REG : REG_GENERIC_NBIT32_6 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => current_PC2_31_port, 
                           DATA_IN(30) => current_PC2_30_port, DATA_IN(29) => 
                           current_PC2_29_port, DATA_IN(28) => 
                           current_PC2_28_port, DATA_IN(27) => 
                           current_PC2_27_port, DATA_IN(26) => 
                           current_PC2_26_port, DATA_IN(25) => 
                           current_PC2_25_port, DATA_IN(24) => 
                           current_PC2_24_port, DATA_IN(23) => 
                           current_PC2_23_port, DATA_IN(22) => 
                           current_PC2_22_port, DATA_IN(21) => 
                           current_PC2_21_port, DATA_IN(20) => 
                           current_PC2_20_port, DATA_IN(19) => 
                           current_PC2_19_port, DATA_IN(18) => 
                           current_PC2_18_port, DATA_IN(17) => 
                           current_PC2_17_port, DATA_IN(16) => 
                           current_PC2_16_port, DATA_IN(15) => 
                           current_PC2_15_port, DATA_IN(14) => 
                           current_PC2_14_port, DATA_IN(13) => 
                           current_PC2_13_port, DATA_IN(12) => 
                           current_PC2_12_port, DATA_IN(11) => 
                           current_PC2_11_port, DATA_IN(10) => 
                           current_PC2_10_port, DATA_IN(9) => 
                           current_PC2_9_port, DATA_IN(8) => current_PC2_8_port
                           , DATA_IN(7) => current_PC2_7_port, DATA_IN(6) => 
                           current_PC2_6_port, DATA_IN(5) => current_PC2_5_port
                           , DATA_IN(4) => current_PC2_4_port, DATA_IN(3) => 
                           current_PC2_3_port, DATA_IN(2) => current_PC2_2_port
                           , DATA_IN(1) => current_PC2_1_port, DATA_IN(0) => 
                           current_PC2_0_port, DATA_OUT(31) => 
                           current_PC3_31_port, DATA_OUT(30) => 
                           current_PC3_30_port, DATA_OUT(29) => 
                           current_PC3_29_port, DATA_OUT(28) => 
                           current_PC3_28_port, DATA_OUT(27) => 
                           current_PC3_27_port, DATA_OUT(26) => 
                           current_PC3_26_port, DATA_OUT(25) => 
                           current_PC3_25_port, DATA_OUT(24) => 
                           current_PC3_24_port, DATA_OUT(23) => 
                           current_PC3_23_port, DATA_OUT(22) => 
                           current_PC3_22_port, DATA_OUT(21) => 
                           current_PC3_21_port, DATA_OUT(20) => 
                           current_PC3_20_port, DATA_OUT(19) => 
                           current_PC3_19_port, DATA_OUT(18) => 
                           current_PC3_18_port, DATA_OUT(17) => 
                           current_PC3_17_port, DATA_OUT(16) => 
                           current_PC3_16_port, DATA_OUT(15) => 
                           current_PC3_15_port, DATA_OUT(14) => 
                           current_PC3_14_port, DATA_OUT(13) => 
                           current_PC3_13_port, DATA_OUT(12) => 
                           current_PC3_12_port, DATA_OUT(11) => 
                           current_PC3_11_port, DATA_OUT(10) => 
                           current_PC3_10_port, DATA_OUT(9) => 
                           current_PC3_9_port, DATA_OUT(8) => 
                           current_PC3_8_port, DATA_OUT(7) => 
                           current_PC3_7_port, DATA_OUT(6) => 
                           current_PC3_6_port, DATA_OUT(5) => 
                           current_PC3_5_port, DATA_OUT(4) => 
                           current_PC3_4_port, DATA_OUT(3) => 
                           current_PC3_3_port, DATA_OUT(2) => 
                           current_PC3_2_port, DATA_OUT(1) => 
                           current_PC3_1_port, DATA_OUT(0) => 
                           current_PC3_0_port);
   NPC_REG : REG_GENERIC_NBIT32_5 port map( CLK => CLK, RST => RST, EN => 
                           NPC_LATCH_EN, DATA_IN(31) => next_NPC_31_port, 
                           DATA_IN(30) => next_NPC_30_port, DATA_IN(29) => 
                           next_NPC_29_port, DATA_IN(28) => next_NPC_28_port, 
                           DATA_IN(27) => next_NPC_27_port, DATA_IN(26) => 
                           next_NPC_26_port, DATA_IN(25) => next_NPC_25_port, 
                           DATA_IN(24) => next_NPC_24_port, DATA_IN(23) => 
                           next_NPC_23_port, DATA_IN(22) => next_NPC_22_port, 
                           DATA_IN(21) => next_NPC_21_port, DATA_IN(20) => 
                           next_NPC_20_port, DATA_IN(19) => next_NPC_19_port, 
                           DATA_IN(18) => next_NPC_18_port, DATA_IN(17) => 
                           next_NPC_17_port, DATA_IN(16) => next_NPC_16_port, 
                           DATA_IN(15) => next_NPC_15_port, DATA_IN(14) => 
                           next_NPC_14_port, DATA_IN(13) => next_NPC_13_port, 
                           DATA_IN(12) => next_NPC_12_port, DATA_IN(11) => 
                           next_NPC_11_port, DATA_IN(10) => next_NPC_10_port, 
                           DATA_IN(9) => next_NPC_9_port, DATA_IN(8) => 
                           next_NPC_8_port, DATA_IN(7) => next_NPC_7_port, 
                           DATA_IN(6) => next_NPC_6_port, DATA_IN(5) => 
                           next_NPC_5_port, DATA_IN(4) => next_NPC_4_port, 
                           DATA_IN(3) => next_NPC_3_port, DATA_IN(2) => 
                           next_NPC_2_port, DATA_IN(1) => next_NPC_1_port, 
                           DATA_IN(0) => next_NPC_0_port, DATA_OUT(31) => 
                           current_NPC_31_port, DATA_OUT(30) => 
                           current_NPC_30_port, DATA_OUT(29) => 
                           current_NPC_29_port, DATA_OUT(28) => 
                           current_NPC_28_port, DATA_OUT(27) => 
                           current_NPC_27_port, DATA_OUT(26) => 
                           current_NPC_26_port, DATA_OUT(25) => 
                           current_NPC_25_port, DATA_OUT(24) => 
                           current_NPC_24_port, DATA_OUT(23) => 
                           current_NPC_23_port, DATA_OUT(22) => 
                           current_NPC_22_port, DATA_OUT(21) => 
                           current_NPC_21_port, DATA_OUT(20) => 
                           current_NPC_20_port, DATA_OUT(19) => 
                           current_NPC_19_port, DATA_OUT(18) => 
                           current_NPC_18_port, DATA_OUT(17) => 
                           current_NPC_17_port, DATA_OUT(16) => 
                           current_NPC_16_port, DATA_OUT(15) => 
                           current_NPC_15_port, DATA_OUT(14) => 
                           current_NPC_14_port, DATA_OUT(13) => 
                           current_NPC_13_port, DATA_OUT(12) => 
                           current_NPC_12_port, DATA_OUT(11) => 
                           current_NPC_11_port, DATA_OUT(10) => 
                           current_NPC_10_port, DATA_OUT(9) => 
                           current_NPC_9_port, DATA_OUT(8) => 
                           current_NPC_8_port, DATA_OUT(7) => 
                           current_NPC_7_port, DATA_OUT(6) => 
                           current_NPC_6_port, DATA_OUT(5) => 
                           current_NPC_5_port, DATA_OUT(4) => 
                           current_NPC_4_port, DATA_OUT(3) => 
                           current_NPC_3_port, DATA_OUT(2) => 
                           current_NPC_2_port, DATA_OUT(1) => 
                           current_NPC_1_port, DATA_OUT(0) => 
                           current_NPC_0_port);
   IR_REG : REG_GENERIC_NBIT32_4 port map( CLK => CLK, RST => RST, EN => 
                           IR_LATCH_EN, DATA_IN(31) => IR_IN(31), DATA_IN(30) 
                           => IR_IN(30), DATA_IN(29) => IR_IN(29), DATA_IN(28) 
                           => IR_IN(28), DATA_IN(27) => IR_IN(27), DATA_IN(26) 
                           => IR_IN(26), DATA_IN(25) => IR_IN(25), DATA_IN(24) 
                           => IR_IN(24), DATA_IN(23) => IR_IN(23), DATA_IN(22) 
                           => IR_IN(22), DATA_IN(21) => IR_IN(21), DATA_IN(20) 
                           => IR_IN(20), DATA_IN(19) => IR_IN(19), DATA_IN(18) 
                           => IR_IN(18), DATA_IN(17) => IR_IN(17), DATA_IN(16) 
                           => IR_IN(16), DATA_IN(15) => IR_IN(15), DATA_IN(14) 
                           => IR_IN(14), DATA_IN(13) => IR_IN(13), DATA_IN(12) 
                           => IR_IN(12), DATA_IN(11) => IR_IN(11), DATA_IN(10) 
                           => IR_IN(10), DATA_IN(9) => IR_IN(9), DATA_IN(8) => 
                           IR_IN(8), DATA_IN(7) => IR_IN(7), DATA_IN(6) => 
                           IR_IN(6), DATA_IN(5) => IR_IN(5), DATA_IN(4) => 
                           IR_IN(4), DATA_IN(3) => IR_IN(3), DATA_IN(2) => 
                           IR_IN(2), DATA_IN(1) => IR_IN(1), DATA_IN(0) => 
                           IR_IN(0), DATA_OUT(31) => n_2386, DATA_OUT(30) => 
                           n_2387, DATA_OUT(29) => n_2388, DATA_OUT(28) => 
                           n_2389, DATA_OUT(27) => n_2390, DATA_OUT(26) => 
                           n_2391, DATA_OUT(25) => current_IW_25_port, 
                           DATA_OUT(24) => current_IW_24_port, DATA_OUT(23) => 
                           current_IW_23_port, DATA_OUT(22) => 
                           current_IW_22_port, DATA_OUT(21) => 
                           current_IW_21_port, DATA_OUT(20) => 
                           current_IW_20_port, DATA_OUT(19) => 
                           current_IW_19_port, DATA_OUT(18) => 
                           current_IW_18_port, DATA_OUT(17) => 
                           current_IW_17_port, DATA_OUT(16) => 
                           current_IW_16_port, DATA_OUT(15) => 
                           current_IW_15_port, DATA_OUT(14) => 
                           current_IW_14_port, DATA_OUT(13) => 
                           current_IW_13_port, DATA_OUT(12) => 
                           current_IW_12_port, DATA_OUT(11) => 
                           current_IW_11_port, DATA_OUT(10) => 
                           current_IW_10_port, DATA_OUT(9) => current_IW_9_port
                           , DATA_OUT(8) => current_IW_8_port, DATA_OUT(7) => 
                           current_IW_7_port, DATA_OUT(6) => current_IW_6_port,
                           DATA_OUT(5) => current_IW_5_port, DATA_OUT(4) => 
                           current_IW_4_port, DATA_OUT(3) => current_IW_3_port,
                           DATA_OUT(2) => current_IW_2_port, DATA_OUT(1) => 
                           current_IW_1_port, DATA_OUT(0) => current_IW_0_port)
                           ;
   IMM_REG : REG_GENERIC_NBIT26 port map( CLK => CLK, RST => RST, EN => 
                           RegIMM_LATCH_EN, DATA_IN(25) => current_IW_25_port, 
                           DATA_IN(24) => current_IW_24_port, DATA_IN(23) => 
                           current_IW_23_port, DATA_IN(22) => 
                           current_IW_22_port, DATA_IN(21) => 
                           current_IW_21_port, DATA_IN(20) => 
                           current_IW_20_port, DATA_IN(19) => 
                           current_IW_19_port, DATA_IN(18) => 
                           current_IW_18_port, DATA_IN(17) => 
                           current_IW_17_port, DATA_IN(16) => 
                           current_IW_16_port, DATA_IN(15) => 
                           current_IW_15_port, DATA_IN(14) => 
                           current_IW_14_port, DATA_IN(13) => 
                           current_IW_13_port, DATA_IN(12) => 
                           current_IW_12_port, DATA_IN(11) => 
                           current_IW_11_port, DATA_IN(10) => 
                           current_IW_10_port, DATA_IN(9) => current_IW_9_port,
                           DATA_IN(8) => current_IW_8_port, DATA_IN(7) => 
                           current_IW_7_port, DATA_IN(6) => current_IW_6_port, 
                           DATA_IN(5) => current_IW_5_port, DATA_IN(4) => 
                           current_IW_4_port, DATA_IN(3) => current_IW_3_port, 
                           DATA_IN(2) => current_IW_2_port, DATA_IN(1) => 
                           current_IW_1_port, DATA_IN(0) => current_IW_0_port, 
                           DATA_OUT(25) => IMM_IN_25_port, DATA_OUT(24) => 
                           IMM_IN_24_port, DATA_OUT(23) => IMM_IN_23_port, 
                           DATA_OUT(22) => IMM_IN_22_port, DATA_OUT(21) => 
                           IMM_IN_21_port, DATA_OUT(20) => IMM_IN_20_port, 
                           DATA_OUT(19) => IMM_IN_19_port, DATA_OUT(18) => 
                           IMM_IN_18_port, DATA_OUT(17) => IMM_IN_17_port, 
                           DATA_OUT(16) => IMM_IN_16_port, DATA_OUT(15) => 
                           IMM_IN_15_port, DATA_OUT(14) => IMM_IN_14_port, 
                           DATA_OUT(13) => IMM_IN_13_port, DATA_OUT(12) => 
                           IMM_IN_12_port, DATA_OUT(11) => IMM_IN_11_port, 
                           DATA_OUT(10) => IMM_IN_10_port, DATA_OUT(9) => 
                           IMM_IN_9_port, DATA_OUT(8) => IMM_IN_8_port, 
                           DATA_OUT(7) => IMM_IN_7_port, DATA_OUT(6) => 
                           IMM_IN_6_port, DATA_OUT(5) => IMM_IN_5_port, 
                           DATA_OUT(4) => IMM_IN_4_port, DATA_OUT(3) => 
                           IMM_IN_3_port, DATA_OUT(2) => IMM_IN_2_port, 
                           DATA_OUT(1) => IMM_IN_1_port, DATA_OUT(0) => 
                           IMM_IN_0_port);
   WB1_REG : REG_GENERIC_NBIT5_0 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, DATA_IN(4) => WB1_IN_4_port, 
                           DATA_IN(3) => WB1_IN_3_port, DATA_IN(2) => 
                           WB1_IN_2_port, DATA_IN(1) => WB1_IN_1_port, 
                           DATA_IN(0) => WB1_IN_0_port, DATA_OUT(4) => 
                           WB2_IN_4_port, DATA_OUT(3) => WB2_IN_3_port, 
                           DATA_OUT(2) => WB2_IN_2_port, DATA_OUT(1) => 
                           WB2_IN_1_port, DATA_OUT(0) => WB2_IN_0_port);
   WB2_REG : REG_GENERIC_NBIT5_2 port map( CLK => CLK, RST => RST, EN => 
                           ALU_OUTREG_EN, DATA_IN(4) => WB2_IN_4_port, 
                           DATA_IN(3) => WB2_IN_3_port, DATA_IN(2) => 
                           WB2_IN_2_port, DATA_IN(1) => WB2_IN_1_port, 
                           DATA_IN(0) => WB2_IN_0_port, DATA_OUT(4) => 
                           WB2_OUT_4_port, DATA_OUT(3) => WB2_OUT_3_port, 
                           DATA_OUT(2) => WB2_OUT_2_port, DATA_OUT(1) => 
                           WB2_OUT_1_port, DATA_OUT(0) => WB2_OUT_0_port);
   WB3_REG : REG_GENERIC_NBIT5_1 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, DATA_IN(4) => WB2_OUT_4_port, 
                           DATA_IN(3) => WB2_OUT_3_port, DATA_IN(2) => 
                           WB2_OUT_2_port, DATA_IN(1) => WB2_OUT_1_port, 
                           DATA_IN(0) => WB2_OUT_0_port, DATA_OUT(4) => 
                           WB3_OUT_4_port, DATA_OUT(3) => WB3_OUT_3_port, 
                           DATA_OUT(2) => WB3_OUT_2_port, DATA_OUT(1) => 
                           WB3_OUT_1_port, DATA_OUT(0) => WB3_OUT_0_port);
   ALU_OUT_REG : REG_GENERIC_NBIT32_3 port map( CLK => CLK, RST => RST, EN => 
                           ALU_OUTREG_EN, DATA_IN(31) => next_ALU_OUT_31_port, 
                           DATA_IN(30) => next_ALU_OUT_30_port, DATA_IN(29) => 
                           next_ALU_OUT_29_port, DATA_IN(28) => 
                           next_ALU_OUT_28_port, DATA_IN(27) => 
                           next_ALU_OUT_27_port, DATA_IN(26) => 
                           next_ALU_OUT_26_port, DATA_IN(25) => 
                           next_ALU_OUT_25_port, DATA_IN(24) => 
                           next_ALU_OUT_24_port, DATA_IN(23) => 
                           next_ALU_OUT_23_port, DATA_IN(22) => 
                           next_ALU_OUT_22_port, DATA_IN(21) => 
                           next_ALU_OUT_21_port, DATA_IN(20) => 
                           next_ALU_OUT_20_port, DATA_IN(19) => 
                           next_ALU_OUT_19_port, DATA_IN(18) => 
                           next_ALU_OUT_18_port, DATA_IN(17) => 
                           next_ALU_OUT_17_port, DATA_IN(16) => 
                           next_ALU_OUT_16_port, DATA_IN(15) => 
                           next_ALU_OUT_15_port, DATA_IN(14) => 
                           next_ALU_OUT_14_port, DATA_IN(13) => 
                           next_ALU_OUT_13_port, DATA_IN(12) => 
                           next_ALU_OUT_12_port, DATA_IN(11) => 
                           next_ALU_OUT_11_port, DATA_IN(10) => 
                           next_ALU_OUT_10_port, DATA_IN(9) => 
                           next_ALU_OUT_9_port, DATA_IN(8) => 
                           next_ALU_OUT_8_port, DATA_IN(7) => 
                           next_ALU_OUT_7_port, DATA_IN(6) => 
                           next_ALU_OUT_6_port, DATA_IN(5) => 
                           next_ALU_OUT_5_port, DATA_IN(4) => 
                           next_ALU_OUT_4_port, DATA_IN(3) => 
                           next_ALU_OUT_3_port, DATA_IN(2) => 
                           next_ALU_OUT_2_port, DATA_IN(1) => 
                           next_ALU_OUT_1_port, DATA_IN(0) => 
                           next_ALU_OUT_0_port, DATA_OUT(31) => 
                           current_ALU_OUT_31_port, DATA_OUT(30) => 
                           current_ALU_OUT_30_port, DATA_OUT(29) => 
                           current_ALU_OUT_29_port, DATA_OUT(28) => 
                           current_ALU_OUT_28_port, DATA_OUT(27) => 
                           current_ALU_OUT_27_port, DATA_OUT(26) => 
                           current_ALU_OUT_26_port, DATA_OUT(25) => 
                           current_ALU_OUT_25_port, DATA_OUT(24) => 
                           current_ALU_OUT_24_port, DATA_OUT(23) => 
                           current_ALU_OUT_23_port, DATA_OUT(22) => 
                           current_ALU_OUT_22_port, DATA_OUT(21) => 
                           current_ALU_OUT_21_port, DATA_OUT(20) => 
                           current_ALU_OUT_20_port, DATA_OUT(19) => 
                           current_ALU_OUT_19_port, DATA_OUT(18) => 
                           current_ALU_OUT_18_port, DATA_OUT(17) => 
                           current_ALU_OUT_17_port, DATA_OUT(16) => 
                           current_ALU_OUT_16_port, DATA_OUT(15) => 
                           current_ALU_OUT_15_port, DATA_OUT(14) => 
                           current_ALU_OUT_14_port, DATA_OUT(13) => 
                           current_ALU_OUT_13_port, DATA_OUT(12) => 
                           current_ALU_OUT_12_port, DATA_OUT(11) => 
                           current_ALU_OUT_11_port, DATA_OUT(10) => 
                           current_ALU_OUT_10_port, DATA_OUT(9) => 
                           current_ALU_OUT_9_port, DATA_OUT(8) => 
                           current_ALU_OUT_8_port, DATA_OUT(7) => 
                           current_ALU_OUT_7_port, DATA_OUT(6) => 
                           current_ALU_OUT_6_port, DATA_OUT(5) => D_ADDR_5_port
                           , DATA_OUT(4) => D_ADDR_4_port, DATA_OUT(3) => 
                           D_ADDR_3_port, DATA_OUT(2) => D_ADDR_2_port, 
                           DATA_OUT(1) => D_ADDR_1_port, DATA_OUT(0) => 
                           D_ADDR_0_port);
   B_OUT_REG : REG_GENERIC_NBIT32_2 port map( CLK => CLK, RST => RST, EN => 
                           ALU_OUTREG_EN, DATA_IN(31) => B_OUT_31_port, 
                           DATA_IN(30) => B_OUT_30_port, DATA_IN(29) => 
                           B_OUT_29_port, DATA_IN(28) => B_OUT_28_port, 
                           DATA_IN(27) => B_OUT_27_port, DATA_IN(26) => 
                           B_OUT_26_port, DATA_IN(25) => B_OUT_25_port, 
                           DATA_IN(24) => B_OUT_24_port, DATA_IN(23) => 
                           B_OUT_23_port, DATA_IN(22) => B_OUT_22_port, 
                           DATA_IN(21) => B_OUT_21_port, DATA_IN(20) => 
                           B_OUT_20_port, DATA_IN(19) => B_OUT_19_port, 
                           DATA_IN(18) => B_OUT_18_port, DATA_IN(17) => 
                           B_OUT_17_port, DATA_IN(16) => B_OUT_16_port, 
                           DATA_IN(15) => B_OUT_15_port, DATA_IN(14) => 
                           B_OUT_14_port, DATA_IN(13) => B_OUT_13_port, 
                           DATA_IN(12) => B_OUT_12_port, DATA_IN(11) => 
                           B_OUT_11_port, DATA_IN(10) => B_OUT_10_port, 
                           DATA_IN(9) => B_OUT_9_port, DATA_IN(8) => 
                           B_OUT_8_port, DATA_IN(7) => B_OUT_7_port, DATA_IN(6)
                           => B_OUT_6_port, DATA_IN(5) => B_OUT_5_port, 
                           DATA_IN(4) => n1, DATA_IN(3) => n2, DATA_IN(2) => 
                           B_OUT_2_port, DATA_IN(1) => n9, DATA_IN(0) => 
                           B_OUT_0_port, DATA_OUT(31) => D_DATA_IN(31), 
                           DATA_OUT(30) => D_DATA_IN(30), DATA_OUT(29) => 
                           D_DATA_IN(29), DATA_OUT(28) => D_DATA_IN(28), 
                           DATA_OUT(27) => D_DATA_IN(27), DATA_OUT(26) => 
                           D_DATA_IN(26), DATA_OUT(25) => D_DATA_IN(25), 
                           DATA_OUT(24) => D_DATA_IN(24), DATA_OUT(23) => 
                           D_DATA_IN(23), DATA_OUT(22) => D_DATA_IN(22), 
                           DATA_OUT(21) => D_DATA_IN(21), DATA_OUT(20) => 
                           D_DATA_IN(20), DATA_OUT(19) => D_DATA_IN(19), 
                           DATA_OUT(18) => D_DATA_IN(18), DATA_OUT(17) => 
                           D_DATA_IN(17), DATA_OUT(16) => D_DATA_IN(16), 
                           DATA_OUT(15) => D_DATA_IN(15), DATA_OUT(14) => 
                           D_DATA_IN(14), DATA_OUT(13) => D_DATA_IN(13), 
                           DATA_OUT(12) => D_DATA_IN(12), DATA_OUT(11) => 
                           D_DATA_IN(11), DATA_OUT(10) => D_DATA_IN(10), 
                           DATA_OUT(9) => D_DATA_IN(9), DATA_OUT(8) => 
                           D_DATA_IN(8), DATA_OUT(7) => D_DATA_IN(7), 
                           DATA_OUT(6) => D_DATA_IN(6), DATA_OUT(5) => 
                           D_DATA_IN(5), DATA_OUT(4) => D_DATA_IN(4), 
                           DATA_OUT(3) => D_DATA_IN(3), DATA_OUT(2) => 
                           D_DATA_IN(2), DATA_OUT(1) => D_DATA_IN(1), 
                           DATA_OUT(0) => D_DATA_IN(0));
   ALU_OUT_REG2 : REG_GENERIC_NBIT32_1 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, DATA_IN(31) => 
                           current_ALU_OUT_31_port, DATA_IN(30) => 
                           current_ALU_OUT_30_port, DATA_IN(29) => 
                           current_ALU_OUT_29_port, DATA_IN(28) => 
                           current_ALU_OUT_28_port, DATA_IN(27) => 
                           current_ALU_OUT_27_port, DATA_IN(26) => 
                           current_ALU_OUT_26_port, DATA_IN(25) => 
                           current_ALU_OUT_25_port, DATA_IN(24) => 
                           current_ALU_OUT_24_port, DATA_IN(23) => 
                           current_ALU_OUT_23_port, DATA_IN(22) => 
                           current_ALU_OUT_22_port, DATA_IN(21) => 
                           current_ALU_OUT_21_port, DATA_IN(20) => 
                           current_ALU_OUT_20_port, DATA_IN(19) => 
                           current_ALU_OUT_19_port, DATA_IN(18) => 
                           current_ALU_OUT_18_port, DATA_IN(17) => 
                           current_ALU_OUT_17_port, DATA_IN(16) => 
                           current_ALU_OUT_16_port, DATA_IN(15) => 
                           current_ALU_OUT_15_port, DATA_IN(14) => 
                           current_ALU_OUT_14_port, DATA_IN(13) => 
                           current_ALU_OUT_13_port, DATA_IN(12) => 
                           current_ALU_OUT_12_port, DATA_IN(11) => 
                           current_ALU_OUT_11_port, DATA_IN(10) => 
                           current_ALU_OUT_10_port, DATA_IN(9) => 
                           current_ALU_OUT_9_port, DATA_IN(8) => 
                           current_ALU_OUT_8_port, DATA_IN(7) => 
                           current_ALU_OUT_7_port, DATA_IN(6) => 
                           current_ALU_OUT_6_port, DATA_IN(5) => n8, DATA_IN(4)
                           => n7, DATA_IN(3) => n6, DATA_IN(2) => n5, 
                           DATA_IN(1) => n4, DATA_IN(0) => n3, DATA_OUT(31) => 
                           current_ALU_OUT2_31_port, DATA_OUT(30) => 
                           current_ALU_OUT2_30_port, DATA_OUT(29) => 
                           current_ALU_OUT2_29_port, DATA_OUT(28) => 
                           current_ALU_OUT2_28_port, DATA_OUT(27) => 
                           current_ALU_OUT2_27_port, DATA_OUT(26) => 
                           current_ALU_OUT2_26_port, DATA_OUT(25) => 
                           current_ALU_OUT2_25_port, DATA_OUT(24) => 
                           current_ALU_OUT2_24_port, DATA_OUT(23) => 
                           current_ALU_OUT2_23_port, DATA_OUT(22) => 
                           current_ALU_OUT2_22_port, DATA_OUT(21) => 
                           current_ALU_OUT2_21_port, DATA_OUT(20) => 
                           current_ALU_OUT2_20_port, DATA_OUT(19) => 
                           current_ALU_OUT2_19_port, DATA_OUT(18) => 
                           current_ALU_OUT2_18_port, DATA_OUT(17) => 
                           current_ALU_OUT2_17_port, DATA_OUT(16) => 
                           current_ALU_OUT2_16_port, DATA_OUT(15) => 
                           current_ALU_OUT2_15_port, DATA_OUT(14) => 
                           current_ALU_OUT2_14_port, DATA_OUT(13) => 
                           current_ALU_OUT2_13_port, DATA_OUT(12) => 
                           current_ALU_OUT2_12_port, DATA_OUT(11) => 
                           current_ALU_OUT2_11_port, DATA_OUT(10) => 
                           current_ALU_OUT2_10_port, DATA_OUT(9) => 
                           current_ALU_OUT2_9_port, DATA_OUT(8) => 
                           current_ALU_OUT2_8_port, DATA_OUT(7) => 
                           current_ALU_OUT2_7_port, DATA_OUT(6) => 
                           current_ALU_OUT2_6_port, DATA_OUT(5) => 
                           current_ALU_OUT2_5_port, DATA_OUT(4) => 
                           current_ALU_OUT2_4_port, DATA_OUT(3) => 
                           current_ALU_OUT2_3_port, DATA_OUT(2) => 
                           current_ALU_OUT2_2_port, DATA_OUT(1) => 
                           current_ALU_OUT2_1_port, DATA_OUT(0) => 
                           current_ALU_OUT2_0_port);
   BU : BRANCHING_UNIT_N32 port map( CLK => CLK, RST => RST, Reg_A(31) => 
                           A_OUT_31_port, Reg_A(30) => A_OUT_30_port, Reg_A(29)
                           => A_OUT_29_port, Reg_A(28) => A_OUT_28_port, 
                           Reg_A(27) => A_OUT_27_port, Reg_A(26) => 
                           A_OUT_26_port, Reg_A(25) => A_OUT_25_port, Reg_A(24)
                           => A_OUT_24_port, Reg_A(23) => A_OUT_23_port, 
                           Reg_A(22) => A_OUT_22_port, Reg_A(21) => 
                           A_OUT_21_port, Reg_A(20) => A_OUT_20_port, Reg_A(19)
                           => A_OUT_19_port, Reg_A(18) => A_OUT_18_port, 
                           Reg_A(17) => A_OUT_17_port, Reg_A(16) => 
                           A_OUT_16_port, Reg_A(15) => A_OUT_15_port, Reg_A(14)
                           => A_OUT_14_port, Reg_A(13) => A_OUT_13_port, 
                           Reg_A(12) => A_OUT_12_port, Reg_A(11) => 
                           A_OUT_11_port, Reg_A(10) => A_OUT_10_port, Reg_A(9) 
                           => A_OUT_9_port, Reg_A(8) => A_OUT_8_port, Reg_A(7) 
                           => A_OUT_7_port, Reg_A(6) => A_OUT_6_port, Reg_A(5) 
                           => A_OUT_5_port, Reg_A(4) => A_OUT_4_port, Reg_A(3) 
                           => A_OUT_3_port, Reg_A(2) => A_OUT_2_port, Reg_A(1) 
                           => A_OUT_1_port, Reg_A(0) => A_OUT_0_port, EQ_cond 
                           => EQ_COND, IS_JUMP => IS_JUMP, branch_taken => 
                           branch_taken);
   PC_MUX : MUX21_GENERIC_NBIT32_0 port map( A(31) => current_NPC_31_port, 
                           A(30) => current_NPC_30_port, A(29) => 
                           current_NPC_29_port, A(28) => current_NPC_28_port, 
                           A(27) => current_NPC_27_port, A(26) => 
                           current_NPC_26_port, A(25) => current_NPC_25_port, 
                           A(24) => current_NPC_24_port, A(23) => 
                           current_NPC_23_port, A(22) => current_NPC_22_port, 
                           A(21) => current_NPC_21_port, A(20) => 
                           current_NPC_20_port, A(19) => current_NPC_19_port, 
                           A(18) => current_NPC_18_port, A(17) => 
                           current_NPC_17_port, A(16) => current_NPC_16_port, 
                           A(15) => current_NPC_15_port, A(14) => 
                           current_NPC_14_port, A(13) => current_NPC_13_port, 
                           A(12) => current_NPC_12_port, A(11) => 
                           current_NPC_11_port, A(10) => current_NPC_10_port, 
                           A(9) => current_NPC_9_port, A(8) => 
                           current_NPC_8_port, A(7) => current_NPC_7_port, A(6)
                           => current_NPC_6_port, A(5) => current_NPC_5_port, 
                           A(4) => current_NPC_4_port, A(3) => 
                           current_NPC_3_port, A(2) => current_NPC_2_port, A(1)
                           => current_NPC_1_port, A(0) => current_NPC_0_port, 
                           B(31) => current_ALU_OUT_31_port, B(30) => 
                           current_ALU_OUT_30_port, B(29) => 
                           current_ALU_OUT_29_port, B(28) => 
                           current_ALU_OUT_28_port, B(27) => 
                           current_ALU_OUT_27_port, B(26) => 
                           current_ALU_OUT_26_port, B(25) => 
                           current_ALU_OUT_25_port, B(24) => 
                           current_ALU_OUT_24_port, B(23) => 
                           current_ALU_OUT_23_port, B(22) => 
                           current_ALU_OUT_22_port, B(21) => 
                           current_ALU_OUT_21_port, B(20) => 
                           current_ALU_OUT_20_port, B(19) => 
                           current_ALU_OUT_19_port, B(18) => 
                           current_ALU_OUT_18_port, B(17) => 
                           current_ALU_OUT_17_port, B(16) => 
                           current_ALU_OUT_16_port, B(15) => 
                           current_ALU_OUT_15_port, B(14) => 
                           current_ALU_OUT_14_port, B(13) => 
                           current_ALU_OUT_13_port, B(12) => 
                           current_ALU_OUT_12_port, B(11) => 
                           current_ALU_OUT_11_port, B(10) => 
                           current_ALU_OUT_10_port, B(9) => 
                           current_ALU_OUT_9_port, B(8) => 
                           current_ALU_OUT_8_port, B(7) => 
                           current_ALU_OUT_7_port, B(6) => 
                           current_ALU_OUT_6_port, B(5) => n8, B(4) => n7, B(3)
                           => n6, B(2) => n5, B(1) => n4, B(0) => n3, SEL => 
                           PC_MUX_SEL, Y(31) => PC_BUS_31_port, Y(30) => 
                           PC_BUS_30_port, Y(29) => PC_BUS_29_port, Y(28) => 
                           PC_BUS_28_port, Y(27) => PC_BUS_27_port, Y(26) => 
                           PC_BUS_26_port, Y(25) => PC_BUS_25_port, Y(24) => 
                           PC_BUS_24_port, Y(23) => PC_BUS_23_port, Y(22) => 
                           PC_BUS_22_port, Y(21) => PC_BUS_21_port, Y(20) => 
                           PC_BUS_20_port, Y(19) => PC_BUS_19_port, Y(18) => 
                           PC_BUS_18_port, Y(17) => PC_BUS_17_port, Y(16) => 
                           PC_BUS_16_port, Y(15) => PC_BUS_15_port, Y(14) => 
                           PC_BUS_14_port, Y(13) => PC_BUS_13_port, Y(12) => 
                           PC_BUS_12_port, Y(11) => PC_BUS_11_port, Y(10) => 
                           PC_BUS_10_port, Y(9) => PC_BUS_9_port, Y(8) => 
                           PC_BUS_8_port, Y(7) => PC_BUS_7_port, Y(6) => 
                           PC_BUS_6_port, Y(5) => PC_BUS_5_port, Y(4) => 
                           PC_BUS_4_port, Y(3) => PC_BUS_3_port, Y(2) => 
                           PC_BUS_2_port, Y(1) => PC_BUS_1_port, Y(0) => 
                           PC_BUS_0_port);
   J_MUX : MUX21 port map( A => X_Logic0_port, B => branch_taken, SEL => 
                           JUMP_EN, Y => PC_MUX_SEL);
   RD_MUX : MUX21_GENERIC_NBIT5_0 port map( A(4) => current_IW_15_port, A(3) =>
                           current_IW_14_port, A(2) => current_IW_13_port, A(1)
                           => current_IW_12_port, A(0) => current_IW_11_port, 
                           B(4) => current_IW_20_port, B(3) => 
                           current_IW_19_port, B(2) => current_IW_18_port, B(1)
                           => current_IW_17_port, B(0) => current_IW_16_port, 
                           SEL => RegIMM_LATCH_EN, Y(4) => WB1_IN_4_port, Y(3) 
                           => WB1_IN_3_port, Y(2) => WB1_IN_2_port, Y(1) => 
                           WB1_IN_1_port, Y(0) => WB1_IN_0_port);
   OP1_MUX : MUX21_GENERIC_NBIT32_4 port map( A(31) => A_OUT_31_port, A(30) => 
                           A_OUT_30_port, A(29) => A_OUT_29_port, A(28) => 
                           A_OUT_28_port, A(27) => A_OUT_27_port, A(26) => 
                           A_OUT_26_port, A(25) => A_OUT_25_port, A(24) => 
                           A_OUT_24_port, A(23) => A_OUT_23_port, A(22) => 
                           A_OUT_22_port, A(21) => A_OUT_21_port, A(20) => 
                           A_OUT_20_port, A(19) => A_OUT_19_port, A(18) => 
                           A_OUT_18_port, A(17) => A_OUT_17_port, A(16) => 
                           A_OUT_16_port, A(15) => A_OUT_15_port, A(14) => 
                           A_OUT_14_port, A(13) => A_OUT_13_port, A(12) => 
                           A_OUT_12_port, A(11) => A_OUT_11_port, A(10) => 
                           A_OUT_10_port, A(9) => A_OUT_9_port, A(8) => 
                           A_OUT_8_port, A(7) => A_OUT_7_port, A(6) => 
                           A_OUT_6_port, A(5) => A_OUT_5_port, A(4) => 
                           A_OUT_4_port, A(3) => A_OUT_3_port, A(2) => 
                           A_OUT_2_port, A(1) => A_OUT_1_port, A(0) => 
                           A_OUT_0_port, B(31) => current_PC1_31_port, B(30) =>
                           current_PC1_30_port, B(29) => current_PC1_29_port, 
                           B(28) => current_PC1_28_port, B(27) => 
                           current_PC1_27_port, B(26) => current_PC1_26_port, 
                           B(25) => current_PC1_25_port, B(24) => 
                           current_PC1_24_port, B(23) => current_PC1_23_port, 
                           B(22) => current_PC1_22_port, B(21) => 
                           current_PC1_21_port, B(20) => current_PC1_20_port, 
                           B(19) => current_PC1_19_port, B(18) => 
                           current_PC1_18_port, B(17) => current_PC1_17_port, 
                           B(16) => current_PC1_16_port, B(15) => 
                           current_PC1_15_port, B(14) => current_PC1_14_port, 
                           B(13) => current_PC1_13_port, B(12) => 
                           current_PC1_12_port, B(11) => current_PC1_11_port, 
                           B(10) => current_PC1_10_port, B(9) => 
                           current_PC1_9_port, B(8) => current_PC1_8_port, B(7)
                           => current_PC1_7_port, B(6) => current_PC1_6_port, 
                           B(5) => current_PC1_5_port, B(4) => 
                           current_PC1_4_port, B(3) => current_PC1_3_port, B(2)
                           => current_PC1_2_port, B(1) => current_PC1_1_port, 
                           B(0) => current_PC1_0_port, SEL => MUXA_SEL, Y(31) 
                           => ALU_OP1_31_port, Y(30) => ALU_OP1_30_port, Y(29) 
                           => ALU_OP1_29_port, Y(28) => ALU_OP1_28_port, Y(27) 
                           => ALU_OP1_27_port, Y(26) => ALU_OP1_26_port, Y(25) 
                           => ALU_OP1_25_port, Y(24) => ALU_OP1_24_port, Y(23) 
                           => ALU_OP1_23_port, Y(22) => ALU_OP1_22_port, Y(21) 
                           => ALU_OP1_21_port, Y(20) => ALU_OP1_20_port, Y(19) 
                           => ALU_OP1_19_port, Y(18) => ALU_OP1_18_port, Y(17) 
                           => ALU_OP1_17_port, Y(16) => ALU_OP1_16_port, Y(15) 
                           => ALU_OP1_15_port, Y(14) => ALU_OP1_14_port, Y(13) 
                           => ALU_OP1_13_port, Y(12) => ALU_OP1_12_port, Y(11) 
                           => ALU_OP1_11_port, Y(10) => ALU_OP1_10_port, Y(9) 
                           => ALU_OP1_9_port, Y(8) => ALU_OP1_8_port, Y(7) => 
                           ALU_OP1_7_port, Y(6) => ALU_OP1_6_port, Y(5) => 
                           ALU_OP1_5_port, Y(4) => ALU_OP1_4_port, Y(3) => 
                           ALU_OP1_3_port, Y(2) => ALU_OP1_2_port, Y(1) => 
                           ALU_OP1_1_port, Y(0) => ALU_OP1_0_port);
   OP2_MUX : MUX21_GENERIC_NBIT32_3 port map( A(31) => B_OUT_31_port, A(30) => 
                           B_OUT_30_port, A(29) => B_OUT_29_port, A(28) => 
                           B_OUT_28_port, A(27) => B_OUT_27_port, A(26) => 
                           B_OUT_26_port, A(25) => B_OUT_25_port, A(24) => 
                           B_OUT_24_port, A(23) => B_OUT_23_port, A(22) => 
                           B_OUT_22_port, A(21) => B_OUT_21_port, A(20) => 
                           B_OUT_20_port, A(19) => B_OUT_19_port, A(18) => 
                           B_OUT_18_port, A(17) => B_OUT_17_port, A(16) => 
                           B_OUT_16_port, A(15) => B_OUT_15_port, A(14) => 
                           B_OUT_14_port, A(13) => B_OUT_13_port, A(12) => 
                           B_OUT_12_port, A(11) => B_OUT_11_port, A(10) => 
                           B_OUT_10_port, A(9) => B_OUT_9_port, A(8) => 
                           B_OUT_8_port, A(7) => B_OUT_7_port, A(6) => 
                           B_OUT_6_port, A(5) => B_OUT_5_port, A(4) => 
                           B_OUT_4_port, A(3) => B_OUT_3_port, A(2) => 
                           B_OUT_2_port, A(1) => B_OUT_1_port, A(0) => 
                           B_OUT_0_port, B(31) => IMM_OUT_31_port, B(30) => 
                           IMM_OUT_30_port, B(29) => IMM_OUT_29_port, B(28) => 
                           IMM_OUT_28_port, B(27) => IMM_OUT_27_port, B(26) => 
                           IMM_OUT_26_port, B(25) => IMM_OUT_25_port, B(24) => 
                           IMM_OUT_24_port, B(23) => IMM_OUT_23_port, B(22) => 
                           IMM_OUT_22_port, B(21) => IMM_OUT_21_port, B(20) => 
                           IMM_OUT_20_port, B(19) => IMM_OUT_19_port, B(18) => 
                           IMM_OUT_18_port, B(17) => IMM_OUT_17_port, B(16) => 
                           IMM_OUT_16_port, B(15) => IMM_OUT_15_port, B(14) => 
                           IMM_OUT_14_port, B(13) => IMM_OUT_13_port, B(12) => 
                           IMM_OUT_12_port, B(11) => IMM_OUT_11_port, B(10) => 
                           IMM_OUT_10_port, B(9) => IMM_OUT_9_port, B(8) => 
                           IMM_OUT_8_port, B(7) => IMM_OUT_7_port, B(6) => 
                           IMM_OUT_6_port, B(5) => IMM_OUT_5_port, B(4) => 
                           IMM_OUT_4_port, B(3) => IMM_OUT_3_port, B(2) => 
                           IMM_OUT_2_port, B(1) => IMM_OUT_1_port, B(0) => 
                           IMM_OUT_0_port, SEL => MUXB_SEL, Y(31) => 
                           ALU_OP2_31_port, Y(30) => ALU_OP2_30_port, Y(29) => 
                           ALU_OP2_29_port, Y(28) => ALU_OP2_28_port, Y(27) => 
                           ALU_OP2_27_port, Y(26) => ALU_OP2_26_port, Y(25) => 
                           ALU_OP2_25_port, Y(24) => ALU_OP2_24_port, Y(23) => 
                           ALU_OP2_23_port, Y(22) => ALU_OP2_22_port, Y(21) => 
                           ALU_OP2_21_port, Y(20) => ALU_OP2_20_port, Y(19) => 
                           ALU_OP2_19_port, Y(18) => ALU_OP2_18_port, Y(17) => 
                           ALU_OP2_17_port, Y(16) => ALU_OP2_16_port, Y(15) => 
                           ALU_OP2_15_port, Y(14) => ALU_OP2_14_port, Y(13) => 
                           ALU_OP2_13_port, Y(12) => ALU_OP2_12_port, Y(11) => 
                           ALU_OP2_11_port, Y(10) => ALU_OP2_10_port, Y(9) => 
                           ALU_OP2_9_port, Y(8) => ALU_OP2_8_port, Y(7) => 
                           ALU_OP2_7_port, Y(6) => ALU_OP2_6_port, Y(5) => 
                           ALU_OP2_5_port, Y(4) => ALU_OP2_4_port, Y(3) => 
                           ALU_OP2_3_port, Y(2) => ALU_OP2_2_port, Y(1) => 
                           ALU_OP2_1_port, Y(0) => ALU_OP2_0_port);
   OUT_MUX : MUX21_GENERIC_NBIT32_2 port map( A(31) => D_DATA_OUT(31), A(30) =>
                           D_DATA_OUT(30), A(29) => D_DATA_OUT(29), A(28) => 
                           D_DATA_OUT(28), A(27) => D_DATA_OUT(27), A(26) => 
                           D_DATA_OUT(26), A(25) => D_DATA_OUT(25), A(24) => 
                           D_DATA_OUT(24), A(23) => D_DATA_OUT(23), A(22) => 
                           D_DATA_OUT(22), A(21) => D_DATA_OUT(21), A(20) => 
                           D_DATA_OUT(20), A(19) => D_DATA_OUT(19), A(18) => 
                           D_DATA_OUT(18), A(17) => D_DATA_OUT(17), A(16) => 
                           D_DATA_OUT(16), A(15) => D_DATA_OUT(15), A(14) => 
                           D_DATA_OUT(14), A(13) => D_DATA_OUT(13), A(12) => 
                           D_DATA_OUT(12), A(11) => D_DATA_OUT(11), A(10) => 
                           D_DATA_OUT(10), A(9) => D_DATA_OUT(9), A(8) => 
                           D_DATA_OUT(8), A(7) => D_DATA_OUT(7), A(6) => 
                           D_DATA_OUT(6), A(5) => D_DATA_OUT(5), A(4) => 
                           D_DATA_OUT(4), A(3) => D_DATA_OUT(3), A(2) => 
                           D_DATA_OUT(2), A(1) => D_DATA_OUT(1), A(0) => 
                           D_DATA_OUT(0), B(31) => current_ALU_OUT2_31_port, 
                           B(30) => current_ALU_OUT2_30_port, B(29) => 
                           current_ALU_OUT2_29_port, B(28) => 
                           current_ALU_OUT2_28_port, B(27) => 
                           current_ALU_OUT2_27_port, B(26) => 
                           current_ALU_OUT2_26_port, B(25) => 
                           current_ALU_OUT2_25_port, B(24) => 
                           current_ALU_OUT2_24_port, B(23) => 
                           current_ALU_OUT2_23_port, B(22) => 
                           current_ALU_OUT2_22_port, B(21) => 
                           current_ALU_OUT2_21_port, B(20) => 
                           current_ALU_OUT2_20_port, B(19) => 
                           current_ALU_OUT2_19_port, B(18) => 
                           current_ALU_OUT2_18_port, B(17) => 
                           current_ALU_OUT2_17_port, B(16) => 
                           current_ALU_OUT2_16_port, B(15) => 
                           current_ALU_OUT2_15_port, B(14) => 
                           current_ALU_OUT2_14_port, B(13) => 
                           current_ALU_OUT2_13_port, B(12) => 
                           current_ALU_OUT2_12_port, B(11) => 
                           current_ALU_OUT2_11_port, B(10) => 
                           current_ALU_OUT2_10_port, B(9) => 
                           current_ALU_OUT2_9_port, B(8) => 
                           current_ALU_OUT2_8_port, B(7) => 
                           current_ALU_OUT2_7_port, B(6) => 
                           current_ALU_OUT2_6_port, B(5) => 
                           current_ALU_OUT2_5_port, B(4) => 
                           current_ALU_OUT2_4_port, B(3) => 
                           current_ALU_OUT2_3_port, B(2) => 
                           current_ALU_OUT2_2_port, B(1) => 
                           current_ALU_OUT2_1_port, B(0) => 
                           current_ALU_OUT2_0_port, SEL => WB_MUX_SEL, Y(31) =>
                           OUT_MUX_DATA_31_port, Y(30) => OUT_MUX_DATA_30_port,
                           Y(29) => OUT_MUX_DATA_29_port, Y(28) => 
                           OUT_MUX_DATA_28_port, Y(27) => OUT_MUX_DATA_27_port,
                           Y(26) => OUT_MUX_DATA_26_port, Y(25) => 
                           OUT_MUX_DATA_25_port, Y(24) => OUT_MUX_DATA_24_port,
                           Y(23) => OUT_MUX_DATA_23_port, Y(22) => 
                           OUT_MUX_DATA_22_port, Y(21) => OUT_MUX_DATA_21_port,
                           Y(20) => OUT_MUX_DATA_20_port, Y(19) => 
                           OUT_MUX_DATA_19_port, Y(18) => OUT_MUX_DATA_18_port,
                           Y(17) => OUT_MUX_DATA_17_port, Y(16) => 
                           OUT_MUX_DATA_16_port, Y(15) => OUT_MUX_DATA_15_port,
                           Y(14) => OUT_MUX_DATA_14_port, Y(13) => 
                           OUT_MUX_DATA_13_port, Y(12) => OUT_MUX_DATA_12_port,
                           Y(11) => OUT_MUX_DATA_11_port, Y(10) => 
                           OUT_MUX_DATA_10_port, Y(9) => OUT_MUX_DATA_9_port, 
                           Y(8) => OUT_MUX_DATA_8_port, Y(7) => 
                           OUT_MUX_DATA_7_port, Y(6) => OUT_MUX_DATA_6_port, 
                           Y(5) => OUT_MUX_DATA_5_port, Y(4) => 
                           OUT_MUX_DATA_4_port, Y(3) => OUT_MUX_DATA_3_port, 
                           Y(2) => OUT_MUX_DATA_2_port, Y(1) => 
                           OUT_MUX_DATA_1_port, Y(0) => OUT_MUX_DATA_0_port);
   JAL_DATA_MUX : MUX21_GENERIC_NBIT32_1 port map( A(31) => 
                           OUT_MUX_DATA_31_port, A(30) => OUT_MUX_DATA_30_port,
                           A(29) => OUT_MUX_DATA_29_port, A(28) => 
                           OUT_MUX_DATA_28_port, A(27) => OUT_MUX_DATA_27_port,
                           A(26) => OUT_MUX_DATA_26_port, A(25) => 
                           OUT_MUX_DATA_25_port, A(24) => OUT_MUX_DATA_24_port,
                           A(23) => OUT_MUX_DATA_23_port, A(22) => 
                           OUT_MUX_DATA_22_port, A(21) => OUT_MUX_DATA_21_port,
                           A(20) => OUT_MUX_DATA_20_port, A(19) => 
                           OUT_MUX_DATA_19_port, A(18) => OUT_MUX_DATA_18_port,
                           A(17) => OUT_MUX_DATA_17_port, A(16) => 
                           OUT_MUX_DATA_16_port, A(15) => OUT_MUX_DATA_15_port,
                           A(14) => OUT_MUX_DATA_14_port, A(13) => 
                           OUT_MUX_DATA_13_port, A(12) => OUT_MUX_DATA_12_port,
                           A(11) => OUT_MUX_DATA_11_port, A(10) => 
                           OUT_MUX_DATA_10_port, A(9) => OUT_MUX_DATA_9_port, 
                           A(8) => OUT_MUX_DATA_8_port, A(7) => 
                           OUT_MUX_DATA_7_port, A(6) => OUT_MUX_DATA_6_port, 
                           A(5) => OUT_MUX_DATA_5_port, A(4) => 
                           OUT_MUX_DATA_4_port, A(3) => OUT_MUX_DATA_3_port, 
                           A(2) => OUT_MUX_DATA_2_port, A(1) => 
                           OUT_MUX_DATA_1_port, A(0) => OUT_MUX_DATA_0_port, 
                           B(31) => current_PC3_31_port, B(30) => 
                           current_PC3_30_port, B(29) => current_PC3_29_port, 
                           B(28) => current_PC3_28_port, B(27) => 
                           current_PC3_27_port, B(26) => current_PC3_26_port, 
                           B(25) => current_PC3_25_port, B(24) => 
                           current_PC3_24_port, B(23) => current_PC3_23_port, 
                           B(22) => current_PC3_22_port, B(21) => 
                           current_PC3_21_port, B(20) => current_PC3_20_port, 
                           B(19) => current_PC3_19_port, B(18) => 
                           current_PC3_18_port, B(17) => current_PC3_17_port, 
                           B(16) => current_PC3_16_port, B(15) => 
                           current_PC3_15_port, B(14) => current_PC3_14_port, 
                           B(13) => current_PC3_13_port, B(12) => 
                           current_PC3_12_port, B(11) => current_PC3_11_port, 
                           B(10) => current_PC3_10_port, B(9) => 
                           current_PC3_9_port, B(8) => current_PC3_8_port, B(7)
                           => current_PC3_7_port, B(6) => current_PC3_6_port, 
                           B(5) => current_PC3_5_port, B(4) => 
                           current_PC3_4_port, B(3) => current_PC3_3_port, B(2)
                           => current_PC3_2_port, B(1) => current_PC3_1_port, 
                           B(0) => current_PC3_0_port, SEL => IS_JAL, Y(31) => 
                           WB_DATA_31_port, Y(30) => WB_DATA_30_port, Y(29) => 
                           WB_DATA_29_port, Y(28) => WB_DATA_28_port, Y(27) => 
                           WB_DATA_27_port, Y(26) => WB_DATA_26_port, Y(25) => 
                           WB_DATA_25_port, Y(24) => WB_DATA_24_port, Y(23) => 
                           WB_DATA_23_port, Y(22) => WB_DATA_22_port, Y(21) => 
                           WB_DATA_21_port, Y(20) => WB_DATA_20_port, Y(19) => 
                           WB_DATA_19_port, Y(18) => WB_DATA_18_port, Y(17) => 
                           WB_DATA_17_port, Y(16) => WB_DATA_16_port, Y(15) => 
                           WB_DATA_15_port, Y(14) => WB_DATA_14_port, Y(13) => 
                           WB_DATA_13_port, Y(12) => WB_DATA_12_port, Y(11) => 
                           WB_DATA_11_port, Y(10) => WB_DATA_10_port, Y(9) => 
                           WB_DATA_9_port, Y(8) => WB_DATA_8_port, Y(7) => 
                           WB_DATA_7_port, Y(6) => WB_DATA_6_port, Y(5) => 
                           WB_DATA_5_port, Y(4) => WB_DATA_4_port, Y(3) => 
                           WB_DATA_3_port, Y(2) => WB_DATA_2_port, Y(1) => 
                           WB_DATA_1_port, Y(0) => WB_DATA_0_port);
   JAL_ADDR_MUX : MUX21_GENERIC_NBIT5_1 port map( A(4) => WB3_OUT_4_port, A(3) 
                           => WB3_OUT_3_port, A(2) => WB3_OUT_2_port, A(1) => 
                           WB3_OUT_1_port, A(0) => WB3_OUT_0_port, B(4) => 
                           X_Logic1_port, B(3) => X_Logic1_port, B(2) => 
                           X_Logic1_port, B(1) => X_Logic1_port, B(0) => 
                           X_Logic1_port, SEL => IS_JAL, Y(4) => WB_ADDR_4_port
                           , Y(3) => WB_ADDR_3_port, Y(2) => WB_ADDR_2_port, 
                           Y(1) => WB_ADDR_1_port, Y(0) => WB_ADDR_0_port);
   PC_ADDER : ADDER_N32 port map( CURR_ADDR(31) => current_PC_31_port, 
                           CURR_ADDR(30) => current_PC_30_port, CURR_ADDR(29) 
                           => current_PC_29_port, CURR_ADDR(28) => 
                           current_PC_28_port, CURR_ADDR(27) => 
                           current_PC_27_port, CURR_ADDR(26) => 
                           current_PC_26_port, CURR_ADDR(25) => 
                           current_PC_25_port, CURR_ADDR(24) => 
                           current_PC_24_port, CURR_ADDR(23) => 
                           current_PC_23_port, CURR_ADDR(22) => 
                           current_PC_22_port, CURR_ADDR(21) => 
                           current_PC_21_port, CURR_ADDR(20) => 
                           current_PC_20_port, CURR_ADDR(19) => 
                           current_PC_19_port, CURR_ADDR(18) => 
                           current_PC_18_port, CURR_ADDR(17) => 
                           current_PC_17_port, CURR_ADDR(16) => 
                           current_PC_16_port, CURR_ADDR(15) => 
                           current_PC_15_port, CURR_ADDR(14) => 
                           current_PC_14_port, CURR_ADDR(13) => 
                           current_PC_13_port, CURR_ADDR(12) => 
                           current_PC_12_port, CURR_ADDR(11) => 
                           current_PC_11_port, CURR_ADDR(10) => 
                           current_PC_10_port, CURR_ADDR(9) => 
                           current_PC_9_port, CURR_ADDR(8) => current_PC_8_port
                           , CURR_ADDR(7) => current_PC_7_port, CURR_ADDR(6) =>
                           current_PC_6_port, CURR_ADDR(5) => current_PC_5_port
                           , CURR_ADDR(4) => current_PC_4_port, CURR_ADDR(3) =>
                           current_PC_3_port, CURR_ADDR(2) => current_PC_2_port
                           , CURR_ADDR(1) => current_PC_1_port, CURR_ADDR(0) =>
                           current_PC_0_port, NEXT_ADDR(31) => next_NPC_31_port
                           , NEXT_ADDR(30) => next_NPC_30_port, NEXT_ADDR(29) 
                           => next_NPC_29_port, NEXT_ADDR(28) => 
                           next_NPC_28_port, NEXT_ADDR(27) => next_NPC_27_port,
                           NEXT_ADDR(26) => next_NPC_26_port, NEXT_ADDR(25) => 
                           next_NPC_25_port, NEXT_ADDR(24) => next_NPC_24_port,
                           NEXT_ADDR(23) => next_NPC_23_port, NEXT_ADDR(22) => 
                           next_NPC_22_port, NEXT_ADDR(21) => next_NPC_21_port,
                           NEXT_ADDR(20) => next_NPC_20_port, NEXT_ADDR(19) => 
                           next_NPC_19_port, NEXT_ADDR(18) => next_NPC_18_port,
                           NEXT_ADDR(17) => next_NPC_17_port, NEXT_ADDR(16) => 
                           next_NPC_16_port, NEXT_ADDR(15) => next_NPC_15_port,
                           NEXT_ADDR(14) => next_NPC_14_port, NEXT_ADDR(13) => 
                           next_NPC_13_port, NEXT_ADDR(12) => next_NPC_12_port,
                           NEXT_ADDR(11) => next_NPC_11_port, NEXT_ADDR(10) => 
                           next_NPC_10_port, NEXT_ADDR(9) => next_NPC_9_port, 
                           NEXT_ADDR(8) => next_NPC_8_port, NEXT_ADDR(7) => 
                           next_NPC_7_port, NEXT_ADDR(6) => next_NPC_6_port, 
                           NEXT_ADDR(5) => next_NPC_5_port, NEXT_ADDR(4) => 
                           next_NPC_4_port, NEXT_ADDR(3) => next_NPC_3_port, 
                           NEXT_ADDR(2) => next_NPC_2_port, NEXT_ADDR(1) => 
                           next_NPC_1_port, NEXT_ADDR(0) => next_NPC_0_port);
   RF : REGISTER_FILE_NBIT32_NREG32 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, RD1 => RegA_LATCH_EN, RD2 => 
                           RegB_LATCH_EN, WR => RF_WE, ADD_WR(4) => 
                           WB_ADDR_4_port, ADD_WR(3) => WB_ADDR_3_port, 
                           ADD_WR(2) => WB_ADDR_2_port, ADD_WR(1) => 
                           WB_ADDR_1_port, ADD_WR(0) => WB_ADDR_0_port, 
                           ADD_RD1(4) => current_IW_25_port, ADD_RD1(3) => 
                           current_IW_24_port, ADD_RD1(2) => current_IW_23_port
                           , ADD_RD1(1) => current_IW_22_port, ADD_RD1(0) => 
                           current_IW_21_port, ADD_RD2(4) => current_IW_20_port
                           , ADD_RD2(3) => current_IW_19_port, ADD_RD2(2) => 
                           current_IW_18_port, ADD_RD2(1) => current_IW_17_port
                           , ADD_RD2(0) => current_IW_16_port, DATAIN(31) => 
                           WB_DATA_31_port, DATAIN(30) => WB_DATA_30_port, 
                           DATAIN(29) => WB_DATA_29_port, DATAIN(28) => 
                           WB_DATA_28_port, DATAIN(27) => WB_DATA_27_port, 
                           DATAIN(26) => WB_DATA_26_port, DATAIN(25) => 
                           WB_DATA_25_port, DATAIN(24) => WB_DATA_24_port, 
                           DATAIN(23) => WB_DATA_23_port, DATAIN(22) => 
                           WB_DATA_22_port, DATAIN(21) => WB_DATA_21_port, 
                           DATAIN(20) => WB_DATA_20_port, DATAIN(19) => 
                           WB_DATA_19_port, DATAIN(18) => WB_DATA_18_port, 
                           DATAIN(17) => WB_DATA_17_port, DATAIN(16) => 
                           WB_DATA_16_port, DATAIN(15) => WB_DATA_15_port, 
                           DATAIN(14) => WB_DATA_14_port, DATAIN(13) => 
                           WB_DATA_13_port, DATAIN(12) => WB_DATA_12_port, 
                           DATAIN(11) => WB_DATA_11_port, DATAIN(10) => 
                           WB_DATA_10_port, DATAIN(9) => WB_DATA_9_port, 
                           DATAIN(8) => WB_DATA_8_port, DATAIN(7) => 
                           WB_DATA_7_port, DATAIN(6) => WB_DATA_6_port, 
                           DATAIN(5) => WB_DATA_5_port, DATAIN(4) => 
                           WB_DATA_4_port, DATAIN(3) => WB_DATA_3_port, 
                           DATAIN(2) => WB_DATA_2_port, DATAIN(1) => 
                           WB_DATA_1_port, DATAIN(0) => WB_DATA_0_port, 
                           OUT1(31) => A_OUT_31_port, OUT1(30) => A_OUT_30_port
                           , OUT1(29) => A_OUT_29_port, OUT1(28) => 
                           A_OUT_28_port, OUT1(27) => A_OUT_27_port, OUT1(26) 
                           => A_OUT_26_port, OUT1(25) => A_OUT_25_port, 
                           OUT1(24) => A_OUT_24_port, OUT1(23) => A_OUT_23_port
                           , OUT1(22) => A_OUT_22_port, OUT1(21) => 
                           A_OUT_21_port, OUT1(20) => A_OUT_20_port, OUT1(19) 
                           => A_OUT_19_port, OUT1(18) => A_OUT_18_port, 
                           OUT1(17) => A_OUT_17_port, OUT1(16) => A_OUT_16_port
                           , OUT1(15) => A_OUT_15_port, OUT1(14) => 
                           A_OUT_14_port, OUT1(13) => A_OUT_13_port, OUT1(12) 
                           => A_OUT_12_port, OUT1(11) => A_OUT_11_port, 
                           OUT1(10) => A_OUT_10_port, OUT1(9) => A_OUT_9_port, 
                           OUT1(8) => A_OUT_8_port, OUT1(7) => A_OUT_7_port, 
                           OUT1(6) => A_OUT_6_port, OUT1(5) => A_OUT_5_port, 
                           OUT1(4) => A_OUT_4_port, OUT1(3) => A_OUT_3_port, 
                           OUT1(2) => A_OUT_2_port, OUT1(1) => A_OUT_1_port, 
                           OUT1(0) => A_OUT_0_port, OUT2(31) => B_OUT_31_port, 
                           OUT2(30) => B_OUT_30_port, OUT2(29) => B_OUT_29_port
                           , OUT2(28) => B_OUT_28_port, OUT2(27) => 
                           B_OUT_27_port, OUT2(26) => B_OUT_26_port, OUT2(25) 
                           => B_OUT_25_port, OUT2(24) => B_OUT_24_port, 
                           OUT2(23) => B_OUT_23_port, OUT2(22) => B_OUT_22_port
                           , OUT2(21) => B_OUT_21_port, OUT2(20) => 
                           B_OUT_20_port, OUT2(19) => B_OUT_19_port, OUT2(18) 
                           => B_OUT_18_port, OUT2(17) => B_OUT_17_port, 
                           OUT2(16) => B_OUT_16_port, OUT2(15) => B_OUT_15_port
                           , OUT2(14) => B_OUT_14_port, OUT2(13) => 
                           B_OUT_13_port, OUT2(12) => B_OUT_12_port, OUT2(11) 
                           => B_OUT_11_port, OUT2(10) => B_OUT_10_port, OUT2(9)
                           => B_OUT_9_port, OUT2(8) => B_OUT_8_port, OUT2(7) =>
                           B_OUT_7_port, OUT2(6) => B_OUT_6_port, OUT2(5) => 
                           B_OUT_5_port, OUT2(4) => B_OUT_4_port, OUT2(3) => 
                           B_OUT_3_port, OUT2(2) => B_OUT_2_port, OUT2(1) => 
                           B_OUT_1_port, OUT2(0) => B_OUT_0_port);
   EXT : EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26 port map( NOT_EXT_IMM(25) => 
                           IMM_IN_25_port, NOT_EXT_IMM(24) => IMM_IN_24_port, 
                           NOT_EXT_IMM(23) => IMM_IN_23_port, NOT_EXT_IMM(22) 
                           => IMM_IN_22_port, NOT_EXT_IMM(21) => IMM_IN_21_port
                           , NOT_EXT_IMM(20) => IMM_IN_20_port, NOT_EXT_IMM(19)
                           => IMM_IN_19_port, NOT_EXT_IMM(18) => IMM_IN_18_port
                           , NOT_EXT_IMM(17) => IMM_IN_17_port, NOT_EXT_IMM(16)
                           => IMM_IN_16_port, NOT_EXT_IMM(15) => IMM_IN_15_port
                           , NOT_EXT_IMM(14) => IMM_IN_14_port, NOT_EXT_IMM(13)
                           => IMM_IN_13_port, NOT_EXT_IMM(12) => IMM_IN_12_port
                           , NOT_EXT_IMM(11) => IMM_IN_11_port, NOT_EXT_IMM(10)
                           => IMM_IN_10_port, NOT_EXT_IMM(9) => IMM_IN_9_port, 
                           NOT_EXT_IMM(8) => IMM_IN_8_port, NOT_EXT_IMM(7) => 
                           IMM_IN_7_port, NOT_EXT_IMM(6) => IMM_IN_6_port, 
                           NOT_EXT_IMM(5) => IMM_IN_5_port, NOT_EXT_IMM(4) => 
                           IMM_IN_4_port, NOT_EXT_IMM(3) => IMM_IN_3_port, 
                           NOT_EXT_IMM(2) => IMM_IN_2_port, NOT_EXT_IMM(1) => 
                           IMM_IN_1_port, NOT_EXT_IMM(0) => IMM_IN_0_port, 
                           SIGNED_IMM => SIGNED_IMM, IS_JUMP => IS_JUMP, 
                           EXT_IMM(31) => IMM_OUT_31_port, EXT_IMM(30) => 
                           IMM_OUT_30_port, EXT_IMM(29) => IMM_OUT_29_port, 
                           EXT_IMM(28) => IMM_OUT_28_port, EXT_IMM(27) => 
                           IMM_OUT_27_port, EXT_IMM(26) => IMM_OUT_26_port, 
                           EXT_IMM(25) => IMM_OUT_25_port, EXT_IMM(24) => 
                           IMM_OUT_24_port, EXT_IMM(23) => IMM_OUT_23_port, 
                           EXT_IMM(22) => IMM_OUT_22_port, EXT_IMM(21) => 
                           IMM_OUT_21_port, EXT_IMM(20) => IMM_OUT_20_port, 
                           EXT_IMM(19) => IMM_OUT_19_port, EXT_IMM(18) => 
                           IMM_OUT_18_port, EXT_IMM(17) => IMM_OUT_17_port, 
                           EXT_IMM(16) => IMM_OUT_16_port, EXT_IMM(15) => 
                           IMM_OUT_15_port, EXT_IMM(14) => IMM_OUT_14_port, 
                           EXT_IMM(13) => IMM_OUT_13_port, EXT_IMM(12) => 
                           IMM_OUT_12_port, EXT_IMM(11) => IMM_OUT_11_port, 
                           EXT_IMM(10) => IMM_OUT_10_port, EXT_IMM(9) => 
                           IMM_OUT_9_port, EXT_IMM(8) => IMM_OUT_8_port, 
                           EXT_IMM(7) => IMM_OUT_7_port, EXT_IMM(6) => 
                           IMM_OUT_6_port, EXT_IMM(5) => IMM_OUT_5_port, 
                           EXT_IMM(4) => IMM_OUT_4_port, EXT_IMM(3) => 
                           IMM_OUT_3_port, EXT_IMM(2) => IMM_OUT_2_port, 
                           EXT_IMM(1) => IMM_OUT_1_port, EXT_IMM(0) => 
                           IMM_OUT_0_port);
   ALU_i : ALU_N32 port map( FUNC(0) => ALU_OPCODE(0), FUNC(1) => ALU_OPCODE(1)
                           , FUNC(2) => ALU_OPCODE(2), FUNC(3) => ALU_OPCODE(3)
                           , DATA1(31) => ALU_OP1_31_port, DATA1(30) => 
                           ALU_OP1_30_port, DATA1(29) => ALU_OP1_29_port, 
                           DATA1(28) => ALU_OP1_28_port, DATA1(27) => 
                           ALU_OP1_27_port, DATA1(26) => ALU_OP1_26_port, 
                           DATA1(25) => ALU_OP1_25_port, DATA1(24) => 
                           ALU_OP1_24_port, DATA1(23) => ALU_OP1_23_port, 
                           DATA1(22) => ALU_OP1_22_port, DATA1(21) => 
                           ALU_OP1_21_port, DATA1(20) => ALU_OP1_20_port, 
                           DATA1(19) => ALU_OP1_19_port, DATA1(18) => 
                           ALU_OP1_18_port, DATA1(17) => ALU_OP1_17_port, 
                           DATA1(16) => ALU_OP1_16_port, DATA1(15) => 
                           ALU_OP1_15_port, DATA1(14) => ALU_OP1_14_port, 
                           DATA1(13) => ALU_OP1_13_port, DATA1(12) => 
                           ALU_OP1_12_port, DATA1(11) => ALU_OP1_11_port, 
                           DATA1(10) => ALU_OP1_10_port, DATA1(9) => 
                           ALU_OP1_9_port, DATA1(8) => ALU_OP1_8_port, DATA1(7)
                           => ALU_OP1_7_port, DATA1(6) => ALU_OP1_6_port, 
                           DATA1(5) => ALU_OP1_5_port, DATA1(4) => 
                           ALU_OP1_4_port, DATA1(3) => ALU_OP1_3_port, DATA1(2)
                           => ALU_OP1_2_port, DATA1(1) => ALU_OP1_1_port, 
                           DATA1(0) => ALU_OP1_0_port, DATA2(31) => 
                           ALU_OP2_31_port, DATA2(30) => ALU_OP2_30_port, 
                           DATA2(29) => ALU_OP2_29_port, DATA2(28) => 
                           ALU_OP2_28_port, DATA2(27) => ALU_OP2_27_port, 
                           DATA2(26) => ALU_OP2_26_port, DATA2(25) => 
                           ALU_OP2_25_port, DATA2(24) => ALU_OP2_24_port, 
                           DATA2(23) => ALU_OP2_23_port, DATA2(22) => 
                           ALU_OP2_22_port, DATA2(21) => ALU_OP2_21_port, 
                           DATA2(20) => ALU_OP2_20_port, DATA2(19) => 
                           ALU_OP2_19_port, DATA2(18) => ALU_OP2_18_port, 
                           DATA2(17) => ALU_OP2_17_port, DATA2(16) => 
                           ALU_OP2_16_port, DATA2(15) => ALU_OP2_15_port, 
                           DATA2(14) => ALU_OP2_14_port, DATA2(13) => 
                           ALU_OP2_13_port, DATA2(12) => ALU_OP2_12_port, 
                           DATA2(11) => ALU_OP2_11_port, DATA2(10) => 
                           ALU_OP2_10_port, DATA2(9) => ALU_OP2_9_port, 
                           DATA2(8) => ALU_OP2_8_port, DATA2(7) => 
                           ALU_OP2_7_port, DATA2(6) => ALU_OP2_6_port, DATA2(5)
                           => ALU_OP2_5_port, DATA2(4) => ALU_OP2_4_port, 
                           DATA2(3) => ALU_OP2_3_port, DATA2(2) => 
                           ALU_OP2_2_port, DATA2(1) => ALU_OP2_1_port, DATA2(0)
                           => ALU_OP2_0_port, OUTALU(31) => 
                           next_ALU_OUT_31_port, OUTALU(30) => 
                           next_ALU_OUT_30_port, OUTALU(29) => 
                           next_ALU_OUT_29_port, OUTALU(28) => 
                           next_ALU_OUT_28_port, OUTALU(27) => 
                           next_ALU_OUT_27_port, OUTALU(26) => 
                           next_ALU_OUT_26_port, OUTALU(25) => 
                           next_ALU_OUT_25_port, OUTALU(24) => 
                           next_ALU_OUT_24_port, OUTALU(23) => 
                           next_ALU_OUT_23_port, OUTALU(22) => 
                           next_ALU_OUT_22_port, OUTALU(21) => 
                           next_ALU_OUT_21_port, OUTALU(20) => 
                           next_ALU_OUT_20_port, OUTALU(19) => 
                           next_ALU_OUT_19_port, OUTALU(18) => 
                           next_ALU_OUT_18_port, OUTALU(17) => 
                           next_ALU_OUT_17_port, OUTALU(16) => 
                           next_ALU_OUT_16_port, OUTALU(15) => 
                           next_ALU_OUT_15_port, OUTALU(14) => 
                           next_ALU_OUT_14_port, OUTALU(13) => 
                           next_ALU_OUT_13_port, OUTALU(12) => 
                           next_ALU_OUT_12_port, OUTALU(11) => 
                           next_ALU_OUT_11_port, OUTALU(10) => 
                           next_ALU_OUT_10_port, OUTALU(9) => 
                           next_ALU_OUT_9_port, OUTALU(8) => 
                           next_ALU_OUT_8_port, OUTALU(7) => 
                           next_ALU_OUT_7_port, OUTALU(6) => 
                           next_ALU_OUT_6_port, OUTALU(5) => 
                           next_ALU_OUT_5_port, OUTALU(4) => 
                           next_ALU_OUT_4_port, OUTALU(3) => 
                           next_ALU_OUT_3_port, OUTALU(2) => 
                           next_ALU_OUT_2_port, OUTALU(1) => 
                           next_ALU_OUT_1_port, OUTALU(0) => 
                           next_ALU_OUT_0_port);

end SYN_STRUCTURE;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_0 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_0;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_0 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76,
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n_2392,
      n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, 
      n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, 
      n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, 
      n_2420, n_2421, n_2422, n_2423 : std_logic;

begin
   DATA_OUT <= ( DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port );
   
   U3 : BUF_X2 port map( A => n106, Z => n71);
   U4 : BUF_X1 port map( A => n1, Z => n69);
   U5 : BUF_X1 port map( A => n1, Z => n68);
   U6 : BUF_X1 port map( A => n1, Z => n70);
   U7 : AND2_X1 port map( A1 => n2, A2 => n74, ZN => n1);
   U8 : INV_X1 port map( A => n3, ZN => n2);
   U9 : INV_X1 port map( A => RST, ZN => n3);
   U42 : CLKBUF_X3 port map( A => n106, Z => n72);
   U43 : CLKBUF_X3 port map( A => n106, Z => n73);
   U44 : OR2_X1 port map( A1 => EN, A2 => n3, ZN => n74);
   U45 : INV_X1 port map( A => n74, ZN => n106);
   U46 : AOI22_X1 port map( A1 => DATA_OUT_0_port, A2 => n71, B1 => DATA_IN(0),
                           B2 => n68, ZN => n75);
   U47 : INV_X1 port map( A => n75, ZN => n139);
   U48 : AOI22_X1 port map( A1 => DATA_OUT_1_port, A2 => n71, B1 => DATA_IN(1),
                           B2 => n68, ZN => n76);
   U49 : INV_X1 port map( A => n76, ZN => n138);
   U50 : AOI22_X1 port map( A1 => DATA_OUT_2_port, A2 => n71, B1 => DATA_IN(2),
                           B2 => n68, ZN => n77);
   U51 : INV_X1 port map( A => n77, ZN => n137);
   U52 : AOI22_X1 port map( A1 => DATA_OUT_3_port, A2 => n71, B1 => DATA_IN(3),
                           B2 => n68, ZN => n78);
   U53 : INV_X1 port map( A => n78, ZN => n136);
   U54 : AOI22_X1 port map( A1 => DATA_OUT_4_port, A2 => n71, B1 => DATA_IN(4),
                           B2 => n68, ZN => n79);
   U55 : INV_X1 port map( A => n79, ZN => n135);
   U56 : AOI22_X1 port map( A1 => DATA_OUT_5_port, A2 => n71, B1 => DATA_IN(5),
                           B2 => n68, ZN => n80);
   U57 : INV_X1 port map( A => n80, ZN => n134);
   U58 : AOI22_X1 port map( A1 => DATA_OUT_6_port, A2 => n71, B1 => DATA_IN(6),
                           B2 => n68, ZN => n81);
   U59 : INV_X1 port map( A => n81, ZN => n133);
   U60 : AOI22_X1 port map( A1 => DATA_OUT_7_port, A2 => n71, B1 => DATA_IN(7),
                           B2 => n68, ZN => n82);
   U61 : INV_X1 port map( A => n82, ZN => n132);
   U62 : AOI22_X1 port map( A1 => DATA_OUT_8_port, A2 => n71, B1 => DATA_IN(8),
                           B2 => n68, ZN => n83);
   U63 : INV_X1 port map( A => n83, ZN => n131);
   U64 : AOI22_X1 port map( A1 => DATA_OUT_9_port, A2 => n71, B1 => DATA_IN(9),
                           B2 => n68, ZN => n84);
   U65 : INV_X1 port map( A => n84, ZN => n130);
   U66 : AOI22_X1 port map( A1 => DATA_OUT_10_port, A2 => n71, B1 => 
                           DATA_IN(10), B2 => n68, ZN => n85);
   U67 : INV_X1 port map( A => n85, ZN => n129);
   U68 : AOI22_X1 port map( A1 => DATA_OUT_11_port, A2 => n71, B1 => 
                           DATA_IN(11), B2 => n68, ZN => n86);
   U69 : INV_X1 port map( A => n86, ZN => n128);
   U70 : AOI22_X1 port map( A1 => DATA_OUT_12_port, A2 => n72, B1 => 
                           DATA_IN(12), B2 => n69, ZN => n87);
   U71 : INV_X1 port map( A => n87, ZN => n127);
   U72 : AOI22_X1 port map( A1 => DATA_OUT_13_port, A2 => n72, B1 => 
                           DATA_IN(13), B2 => n69, ZN => n88);
   U73 : INV_X1 port map( A => n88, ZN => n126);
   U74 : AOI22_X1 port map( A1 => DATA_OUT_14_port, A2 => n72, B1 => 
                           DATA_IN(14), B2 => n69, ZN => n89);
   U75 : INV_X1 port map( A => n89, ZN => n125);
   U76 : AOI22_X1 port map( A1 => DATA_OUT_15_port, A2 => n72, B1 => 
                           DATA_IN(15), B2 => n69, ZN => n90);
   U77 : INV_X1 port map( A => n90, ZN => n124);
   U78 : AOI22_X1 port map( A1 => DATA_OUT_16_port, A2 => n72, B1 => 
                           DATA_IN(16), B2 => n69, ZN => n91);
   U79 : INV_X1 port map( A => n91, ZN => n123);
   U80 : AOI22_X1 port map( A1 => DATA_OUT_17_port, A2 => n72, B1 => 
                           DATA_IN(17), B2 => n69, ZN => n92);
   U81 : INV_X1 port map( A => n92, ZN => n122);
   U82 : AOI22_X1 port map( A1 => DATA_OUT_18_port, A2 => n72, B1 => 
                           DATA_IN(18), B2 => n69, ZN => n93);
   U83 : INV_X1 port map( A => n93, ZN => n121);
   U84 : AOI22_X1 port map( A1 => DATA_OUT_19_port, A2 => n72, B1 => 
                           DATA_IN(19), B2 => n69, ZN => n94);
   U85 : INV_X1 port map( A => n94, ZN => n120);
   U86 : AOI22_X1 port map( A1 => DATA_OUT_20_port, A2 => n72, B1 => 
                           DATA_IN(20), B2 => n69, ZN => n95);
   U87 : INV_X1 port map( A => n95, ZN => n119);
   U88 : AOI22_X1 port map( A1 => DATA_OUT_21_port, A2 => n72, B1 => 
                           DATA_IN(21), B2 => n69, ZN => n96);
   U89 : INV_X1 port map( A => n96, ZN => n118);
   U90 : AOI22_X1 port map( A1 => DATA_OUT_22_port, A2 => n72, B1 => 
                           DATA_IN(22), B2 => n69, ZN => n97);
   U91 : INV_X1 port map( A => n97, ZN => n117);
   U92 : AOI22_X1 port map( A1 => DATA_OUT_23_port, A2 => n72, B1 => 
                           DATA_IN(23), B2 => n69, ZN => n98);
   U93 : INV_X1 port map( A => n98, ZN => n116);
   U94 : AOI22_X1 port map( A1 => DATA_OUT_24_port, A2 => n73, B1 => 
                           DATA_IN(24), B2 => n70, ZN => n99);
   U95 : INV_X1 port map( A => n99, ZN => n115);
   U96 : AOI22_X1 port map( A1 => DATA_OUT_25_port, A2 => n73, B1 => 
                           DATA_IN(25), B2 => n70, ZN => n100);
   U97 : INV_X1 port map( A => n100, ZN => n114);
   U98 : AOI22_X1 port map( A1 => DATA_OUT_26_port, A2 => n73, B1 => 
                           DATA_IN(26), B2 => n70, ZN => n101);
   U99 : INV_X1 port map( A => n101, ZN => n113);
   U100 : AOI22_X1 port map( A1 => DATA_OUT_27_port, A2 => n73, B1 => 
                           DATA_IN(27), B2 => n70, ZN => n102);
   U101 : INV_X1 port map( A => n102, ZN => n112);
   U102 : AOI22_X1 port map( A1 => DATA_OUT_28_port, A2 => n73, B1 => 
                           DATA_IN(28), B2 => n70, ZN => n103);
   U103 : INV_X1 port map( A => n103, ZN => n111);
   U104 : AOI22_X1 port map( A1 => DATA_OUT_29_port, A2 => n73, B1 => 
                           DATA_IN(29), B2 => n70, ZN => n104);
   U105 : INV_X1 port map( A => n104, ZN => n110);
   U106 : AOI22_X1 port map( A1 => DATA_OUT_30_port, A2 => n73, B1 => 
                           DATA_IN(30), B2 => n70, ZN => n105);
   U107 : INV_X1 port map( A => n105, ZN => n109);
   U108 : AOI22_X1 port map( A1 => DATA_OUT_31_port, A2 => n73, B1 => 
                           DATA_IN(31), B2 => n70, ZN => n107);
   U109 : INV_X1 port map( A => n107, ZN => n108);
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n108, CK => CLK, Q => 
                           DATA_OUT_31_port, QN => n_2392);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n109, CK => CLK, Q => 
                           DATA_OUT_30_port, QN => n_2393);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n110, CK => CLK, Q => 
                           DATA_OUT_29_port, QN => n_2394);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n111, CK => CLK, Q => 
                           DATA_OUT_28_port, QN => n_2395);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n112, CK => CLK, Q => 
                           DATA_OUT_27_port, QN => n_2396);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n113, CK => CLK, Q => 
                           DATA_OUT_26_port, QN => n_2397);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n114, CK => CLK, Q => 
                           DATA_OUT_25_port, QN => n_2398);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n115, CK => CLK, Q => 
                           DATA_OUT_24_port, QN => n_2399);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n128, CK => CLK, Q => 
                           DATA_OUT_11_port, QN => n_2400);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n129, CK => CLK, Q => 
                           DATA_OUT_10_port, QN => n_2401);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n130, CK => CLK, Q => 
                           DATA_OUT_9_port, QN => n_2402);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n131, CK => CLK, Q => 
                           DATA_OUT_8_port, QN => n_2403);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n132, CK => CLK, Q => 
                           DATA_OUT_7_port, QN => n_2404);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n133, CK => CLK, Q => 
                           DATA_OUT_6_port, QN => n_2405);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n134, CK => CLK, Q => 
                           DATA_OUT_5_port, QN => n_2406);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n135, CK => CLK, Q => 
                           DATA_OUT_4_port, QN => n_2407);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n136, CK => CLK, Q => 
                           DATA_OUT_3_port, QN => n_2408);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n137, CK => CLK, Q => 
                           DATA_OUT_2_port, QN => n_2409);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n138, CK => CLK, Q => 
                           DATA_OUT_1_port, QN => n_2410);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n139, CK => CLK, Q => 
                           DATA_OUT_0_port, QN => n_2411);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n116, CK => CLK, Q => 
                           DATA_OUT_23_port, QN => n_2412);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n117, CK => CLK, Q => 
                           DATA_OUT_22_port, QN => n_2413);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n118, CK => CLK, Q => 
                           DATA_OUT_21_port, QN => n_2414);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n119, CK => CLK, Q => 
                           DATA_OUT_20_port, QN => n_2415);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n120, CK => CLK, Q => 
                           DATA_OUT_19_port, QN => n_2416);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n121, CK => CLK, Q => 
                           DATA_OUT_18_port, QN => n_2417);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n122, CK => CLK, Q => 
                           DATA_OUT_17_port, QN => n_2418);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n123, CK => CLK, Q => 
                           DATA_OUT_16_port, QN => n_2419);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n124, CK => CLK, Q => 
                           DATA_OUT_15_port, QN => n_2420);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n125, CK => CLK, Q => 
                           DATA_OUT_14_port, QN => n_2421);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n126, CK => CLK, Q => 
                           DATA_OUT_13_port, QN => n_2422);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n127, CK => CLK, Q => 
                           DATA_OUT_12_port, QN => n_2423);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( CLK, RST : in std_logic;  I_ADDR : out std_logic_vector (31 downto 0);
         I_DATA : in std_logic_vector (31 downto 0);  D_RR, D_WR : out 
         std_logic;  D_ADDR : out std_logic_vector (5 downto 0);  D_DATA_IN : 
         out std_logic_vector (31 downto 0);  D_DATA_OUT : in std_logic_vector 
         (31 downto 0));

end DLX;

architecture SYN_DLX_RTL of DLX is

   component dlx_cu
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
            EQ_COND, IS_JUMP : out std_logic;  ALU_OPCODE : out 
            std_logic_vector (0 to 3);  DRAM_WE, LMD_LATCH_EN, JUMP_EN, 
            PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE : out std_logic);
   end component;
   
   component DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64
      port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
            EQ_COND, IS_JUMP : in std_logic;  ALU_OPCODE : in std_logic_vector 
            (0 to 3);  JUMP_EN, PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE : in 
            std_logic;  D_ADDR : out std_logic_vector (5 downto 0);  D_DATA_IN 
            : out std_logic_vector (31 downto 0);  D_DATA_OUT, PC_IN : in 
            std_logic_vector (31 downto 0);  PC_BUS : out std_logic_vector (31 
            downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_0
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal I_ADDR_31_port, I_ADDR_30_port, I_ADDR_29_port, I_ADDR_28_port, 
      I_ADDR_27_port, I_ADDR_26_port, I_ADDR_25_port, I_ADDR_24_port, 
      I_ADDR_23_port, I_ADDR_22_port, I_ADDR_21_port, I_ADDR_20_port, 
      I_ADDR_19_port, I_ADDR_18_port, I_ADDR_17_port, I_ADDR_16_port, 
      I_ADDR_15_port, I_ADDR_14_port, I_ADDR_13_port, I_ADDR_12_port, 
      I_ADDR_11_port, I_ADDR_10_port, I_ADDR_9_port, I_ADDR_8_port, 
      I_ADDR_7_port, I_ADDR_6_port, I_ADDR_5_port, I_ADDR_4_port, I_ADDR_3_port
      , I_ADDR_2_port, I_ADDR_1_port, I_ADDR_0_port, PC_LATCH_EN, 
      PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, IR_LATCH_EN, NPC_LATCH_EN,
      RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, 
      MUXB_SEL, ALU_OUTREG_EN, EQ_COND, IS_JUMP, ALU_OPCODE_3_port, 
      ALU_OPCODE_2_port, ALU_OPCODE_1_port, ALU_OPCODE_0_port, JUMP_EN, IS_JAL,
      WB_MUX_SEL, RF_WE, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, 
      n28, n29, n30, n31, n32, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, 
      n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, 
      n_2439, n_2440, n_2441 : std_logic;

begin
   I_ADDR <= ( I_ADDR_31_port, I_ADDR_30_port, I_ADDR_29_port, I_ADDR_28_port, 
      I_ADDR_27_port, I_ADDR_26_port, I_ADDR_25_port, I_ADDR_24_port, 
      I_ADDR_23_port, I_ADDR_22_port, I_ADDR_21_port, I_ADDR_20_port, 
      I_ADDR_19_port, I_ADDR_18_port, I_ADDR_17_port, I_ADDR_16_port, 
      I_ADDR_15_port, I_ADDR_14_port, I_ADDR_13_port, I_ADDR_12_port, 
      I_ADDR_11_port, I_ADDR_10_port, I_ADDR_9_port, I_ADDR_8_port, 
      I_ADDR_7_port, I_ADDR_6_port, I_ADDR_5_port, I_ADDR_4_port, I_ADDR_3_port
      , I_ADDR_2_port, I_ADDR_1_port, I_ADDR_0_port );
   
   U1 : CLKBUF_X1 port map( A => I_ADDR_0_port, Z => n1);
   U2 : CLKBUF_X1 port map( A => I_ADDR_1_port, Z => n2);
   U3 : CLKBUF_X1 port map( A => I_ADDR_2_port, Z => n3);
   U4 : CLKBUF_X1 port map( A => I_ADDR_3_port, Z => n4);
   U5 : CLKBUF_X1 port map( A => I_ADDR_4_port, Z => n5);
   U6 : CLKBUF_X1 port map( A => I_ADDR_5_port, Z => n6);
   U7 : CLKBUF_X1 port map( A => I_ADDR_6_port, Z => n7);
   U8 : CLKBUF_X1 port map( A => I_ADDR_7_port, Z => n8);
   U9 : CLKBUF_X1 port map( A => I_ADDR_8_port, Z => n9);
   U10 : CLKBUF_X1 port map( A => I_ADDR_9_port, Z => n10);
   U11 : CLKBUF_X1 port map( A => I_ADDR_10_port, Z => n11);
   U12 : CLKBUF_X1 port map( A => I_ADDR_11_port, Z => n12);
   U13 : CLKBUF_X1 port map( A => I_ADDR_12_port, Z => n13);
   U14 : CLKBUF_X1 port map( A => I_ADDR_13_port, Z => n14);
   U15 : CLKBUF_X1 port map( A => I_ADDR_14_port, Z => n15);
   U16 : CLKBUF_X1 port map( A => I_ADDR_15_port, Z => n16);
   U17 : CLKBUF_X1 port map( A => I_ADDR_16_port, Z => n17);
   U18 : CLKBUF_X1 port map( A => I_ADDR_17_port, Z => n18);
   U19 : CLKBUF_X1 port map( A => I_ADDR_18_port, Z => n19);
   U20 : CLKBUF_X1 port map( A => I_ADDR_19_port, Z => n20);
   U21 : CLKBUF_X1 port map( A => I_ADDR_20_port, Z => n21);
   U22 : CLKBUF_X1 port map( A => I_ADDR_21_port, Z => n22);
   U23 : CLKBUF_X1 port map( A => I_ADDR_22_port, Z => n23);
   U24 : CLKBUF_X1 port map( A => I_ADDR_23_port, Z => n24);
   U25 : CLKBUF_X1 port map( A => I_ADDR_24_port, Z => n25);
   U26 : CLKBUF_X1 port map( A => I_ADDR_25_port, Z => n26);
   U27 : CLKBUF_X1 port map( A => I_ADDR_26_port, Z => n27);
   U28 : CLKBUF_X1 port map( A => I_ADDR_27_port, Z => n28);
   U29 : CLKBUF_X1 port map( A => I_ADDR_28_port, Z => n29);
   U30 : CLKBUF_X1 port map( A => I_ADDR_29_port, Z => n30);
   U31 : CLKBUF_X1 port map( A => I_ADDR_30_port, Z => n31);
   U32 : CLKBUF_X1 port map( A => I_ADDR_31_port, Z => n32);
   RF_WE <= '0';
   WB_MUX_SEL <= '0';
   IS_JAL <= '0';
   PC_LATCH_EN <= '0';
   JUMP_EN <= '0';
   D_RR <= '0';
   D_WR <= '0';
   IS_JUMP <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   SIGNED_IMM <= '0';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   NPC_LATCH_EN <= '0';
   IR_LATCH_EN <= '0';
   PC_REG : REG_GENERIC_NBIT32_0 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => PC_BUS_31_port, 
                           DATA_IN(30) => PC_BUS_30_port, DATA_IN(29) => 
                           PC_BUS_29_port, DATA_IN(28) => PC_BUS_28_port, 
                           DATA_IN(27) => PC_BUS_27_port, DATA_IN(26) => 
                           PC_BUS_26_port, DATA_IN(25) => PC_BUS_25_port, 
                           DATA_IN(24) => PC_BUS_24_port, DATA_IN(23) => 
                           PC_BUS_23_port, DATA_IN(22) => PC_BUS_22_port, 
                           DATA_IN(21) => PC_BUS_21_port, DATA_IN(20) => 
                           PC_BUS_20_port, DATA_IN(19) => PC_BUS_19_port, 
                           DATA_IN(18) => PC_BUS_18_port, DATA_IN(17) => 
                           PC_BUS_17_port, DATA_IN(16) => PC_BUS_16_port, 
                           DATA_IN(15) => PC_BUS_15_port, DATA_IN(14) => 
                           PC_BUS_14_port, DATA_IN(13) => PC_BUS_13_port, 
                           DATA_IN(12) => PC_BUS_12_port, DATA_IN(11) => 
                           PC_BUS_11_port, DATA_IN(10) => PC_BUS_10_port, 
                           DATA_IN(9) => PC_BUS_9_port, DATA_IN(8) => 
                           PC_BUS_8_port, DATA_IN(7) => PC_BUS_7_port, 
                           DATA_IN(6) => PC_BUS_6_port, DATA_IN(5) => 
                           PC_BUS_5_port, DATA_IN(4) => PC_BUS_4_port, 
                           DATA_IN(3) => PC_BUS_3_port, DATA_IN(2) => 
                           PC_BUS_2_port, DATA_IN(1) => PC_BUS_1_port, 
                           DATA_IN(0) => PC_BUS_0_port, DATA_OUT(31) => 
                           I_ADDR_31_port, DATA_OUT(30) => I_ADDR_30_port, 
                           DATA_OUT(29) => I_ADDR_29_port, DATA_OUT(28) => 
                           I_ADDR_28_port, DATA_OUT(27) => I_ADDR_27_port, 
                           DATA_OUT(26) => I_ADDR_26_port, DATA_OUT(25) => 
                           I_ADDR_25_port, DATA_OUT(24) => I_ADDR_24_port, 
                           DATA_OUT(23) => I_ADDR_23_port, DATA_OUT(22) => 
                           I_ADDR_22_port, DATA_OUT(21) => I_ADDR_21_port, 
                           DATA_OUT(20) => I_ADDR_20_port, DATA_OUT(19) => 
                           I_ADDR_19_port, DATA_OUT(18) => I_ADDR_18_port, 
                           DATA_OUT(17) => I_ADDR_17_port, DATA_OUT(16) => 
                           I_ADDR_16_port, DATA_OUT(15) => I_ADDR_15_port, 
                           DATA_OUT(14) => I_ADDR_14_port, DATA_OUT(13) => 
                           I_ADDR_13_port, DATA_OUT(12) => I_ADDR_12_port, 
                           DATA_OUT(11) => I_ADDR_11_port, DATA_OUT(10) => 
                           I_ADDR_10_port, DATA_OUT(9) => I_ADDR_9_port, 
                           DATA_OUT(8) => I_ADDR_8_port, DATA_OUT(7) => 
                           I_ADDR_7_port, DATA_OUT(6) => I_ADDR_6_port, 
                           DATA_OUT(5) => I_ADDR_5_port, DATA_OUT(4) => 
                           I_ADDR_4_port, DATA_OUT(3) => I_ADDR_3_port, 
                           DATA_OUT(2) => I_ADDR_2_port, DATA_OUT(1) => 
                           I_ADDR_1_port, DATA_OUT(0) => I_ADDR_0_port);
   DP : DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 port map( CLK => CLK
                           , RST => RST, IR_IN(31) => I_DATA(31), IR_IN(30) => 
                           I_DATA(30), IR_IN(29) => I_DATA(29), IR_IN(28) => 
                           I_DATA(28), IR_IN(27) => I_DATA(27), IR_IN(26) => 
                           I_DATA(26), IR_IN(25) => I_DATA(25), IR_IN(24) => 
                           I_DATA(24), IR_IN(23) => I_DATA(23), IR_IN(22) => 
                           I_DATA(22), IR_IN(21) => I_DATA(21), IR_IN(20) => 
                           I_DATA(20), IR_IN(19) => I_DATA(19), IR_IN(18) => 
                           I_DATA(18), IR_IN(17) => I_DATA(17), IR_IN(16) => 
                           I_DATA(16), IR_IN(15) => I_DATA(15), IR_IN(14) => 
                           I_DATA(14), IR_IN(13) => I_DATA(13), IR_IN(12) => 
                           I_DATA(12), IR_IN(11) => I_DATA(11), IR_IN(10) => 
                           I_DATA(10), IR_IN(9) => I_DATA(9), IR_IN(8) => 
                           I_DATA(8), IR_IN(7) => I_DATA(7), IR_IN(6) => 
                           I_DATA(6), IR_IN(5) => I_DATA(5), IR_IN(4) => 
                           I_DATA(4), IR_IN(3) => I_DATA(3), IR_IN(2) => 
                           I_DATA(2), IR_IN(1) => I_DATA(1), IR_IN(0) => 
                           I_DATA(0), IR_LATCH_EN => IR_LATCH_EN, NPC_LATCH_EN 
                           => NPC_LATCH_EN, RegA_LATCH_EN => RegA_LATCH_EN, 
                           RegB_LATCH_EN => RegB_LATCH_EN, RegIMM_LATCH_EN => 
                           RegIMM_LATCH_EN, SIGNED_IMM => SIGNED_IMM, MUXA_SEL 
                           => MUXA_SEL, MUXB_SEL => MUXB_SEL, ALU_OUTREG_EN => 
                           ALU_OUTREG_EN, EQ_COND => EQ_COND, IS_JUMP => 
                           IS_JUMP, ALU_OPCODE(0) => ALU_OPCODE_3_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_2_port, ALU_OPCODE(2) =>
                           ALU_OPCODE_1_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_0_port, JUMP_EN => JUMP_EN, PC_LATCH_EN 
                           => PC_LATCH_EN, IS_JAL => IS_JAL, WB_MUX_SEL => 
                           WB_MUX_SEL, RF_WE => RF_WE, D_ADDR(5) => D_ADDR(5), 
                           D_ADDR(4) => D_ADDR(4), D_ADDR(3) => D_ADDR(3), 
                           D_ADDR(2) => D_ADDR(2), D_ADDR(1) => D_ADDR(1), 
                           D_ADDR(0) => D_ADDR(0), D_DATA_IN(31) => 
                           D_DATA_IN(31), D_DATA_IN(30) => D_DATA_IN(30), 
                           D_DATA_IN(29) => D_DATA_IN(29), D_DATA_IN(28) => 
                           D_DATA_IN(28), D_DATA_IN(27) => D_DATA_IN(27), 
                           D_DATA_IN(26) => D_DATA_IN(26), D_DATA_IN(25) => 
                           D_DATA_IN(25), D_DATA_IN(24) => D_DATA_IN(24), 
                           D_DATA_IN(23) => D_DATA_IN(23), D_DATA_IN(22) => 
                           D_DATA_IN(22), D_DATA_IN(21) => D_DATA_IN(21), 
                           D_DATA_IN(20) => D_DATA_IN(20), D_DATA_IN(19) => 
                           D_DATA_IN(19), D_DATA_IN(18) => D_DATA_IN(18), 
                           D_DATA_IN(17) => D_DATA_IN(17), D_DATA_IN(16) => 
                           D_DATA_IN(16), D_DATA_IN(15) => D_DATA_IN(15), 
                           D_DATA_IN(14) => D_DATA_IN(14), D_DATA_IN(13) => 
                           D_DATA_IN(13), D_DATA_IN(12) => D_DATA_IN(12), 
                           D_DATA_IN(11) => D_DATA_IN(11), D_DATA_IN(10) => 
                           D_DATA_IN(10), D_DATA_IN(9) => D_DATA_IN(9), 
                           D_DATA_IN(8) => D_DATA_IN(8), D_DATA_IN(7) => 
                           D_DATA_IN(7), D_DATA_IN(6) => D_DATA_IN(6), 
                           D_DATA_IN(5) => D_DATA_IN(5), D_DATA_IN(4) => 
                           D_DATA_IN(4), D_DATA_IN(3) => D_DATA_IN(3), 
                           D_DATA_IN(2) => D_DATA_IN(2), D_DATA_IN(1) => 
                           D_DATA_IN(1), D_DATA_IN(0) => D_DATA_IN(0), 
                           D_DATA_OUT(31) => D_DATA_OUT(31), D_DATA_OUT(30) => 
                           D_DATA_OUT(30), D_DATA_OUT(29) => D_DATA_OUT(29), 
                           D_DATA_OUT(28) => D_DATA_OUT(28), D_DATA_OUT(27) => 
                           D_DATA_OUT(27), D_DATA_OUT(26) => D_DATA_OUT(26), 
                           D_DATA_OUT(25) => D_DATA_OUT(25), D_DATA_OUT(24) => 
                           D_DATA_OUT(24), D_DATA_OUT(23) => D_DATA_OUT(23), 
                           D_DATA_OUT(22) => D_DATA_OUT(22), D_DATA_OUT(21) => 
                           D_DATA_OUT(21), D_DATA_OUT(20) => D_DATA_OUT(20), 
                           D_DATA_OUT(19) => D_DATA_OUT(19), D_DATA_OUT(18) => 
                           D_DATA_OUT(18), D_DATA_OUT(17) => D_DATA_OUT(17), 
                           D_DATA_OUT(16) => D_DATA_OUT(16), D_DATA_OUT(15) => 
                           D_DATA_OUT(15), D_DATA_OUT(14) => D_DATA_OUT(14), 
                           D_DATA_OUT(13) => D_DATA_OUT(13), D_DATA_OUT(12) => 
                           D_DATA_OUT(12), D_DATA_OUT(11) => D_DATA_OUT(11), 
                           D_DATA_OUT(10) => D_DATA_OUT(10), D_DATA_OUT(9) => 
                           D_DATA_OUT(9), D_DATA_OUT(8) => D_DATA_OUT(8), 
                           D_DATA_OUT(7) => D_DATA_OUT(7), D_DATA_OUT(6) => 
                           D_DATA_OUT(6), D_DATA_OUT(5) => D_DATA_OUT(5), 
                           D_DATA_OUT(4) => D_DATA_OUT(4), D_DATA_OUT(3) => 
                           D_DATA_OUT(3), D_DATA_OUT(2) => D_DATA_OUT(2), 
                           D_DATA_OUT(1) => D_DATA_OUT(1), D_DATA_OUT(0) => 
                           D_DATA_OUT(0), PC_IN(31) => n32, PC_IN(30) => n31, 
                           PC_IN(29) => n30, PC_IN(28) => n29, PC_IN(27) => n28
                           , PC_IN(26) => n27, PC_IN(25) => n26, PC_IN(24) => 
                           n25, PC_IN(23) => n24, PC_IN(22) => n23, PC_IN(21) 
                           => n22, PC_IN(20) => n21, PC_IN(19) => n20, 
                           PC_IN(18) => n19, PC_IN(17) => n18, PC_IN(16) => n17
                           , PC_IN(15) => n16, PC_IN(14) => n15, PC_IN(13) => 
                           n14, PC_IN(12) => n13, PC_IN(11) => n12, PC_IN(10) 
                           => n11, PC_IN(9) => n10, PC_IN(8) => n9, PC_IN(7) =>
                           n8, PC_IN(6) => n7, PC_IN(5) => n6, PC_IN(4) => n5, 
                           PC_IN(3) => n4, PC_IN(2) => n3, PC_IN(1) => n2, 
                           PC_IN(0) => n1, PC_BUS(31) => PC_BUS_31_port, 
                           PC_BUS(30) => PC_BUS_30_port, PC_BUS(29) => 
                           PC_BUS_29_port, PC_BUS(28) => PC_BUS_28_port, 
                           PC_BUS(27) => PC_BUS_27_port, PC_BUS(26) => 
                           PC_BUS_26_port, PC_BUS(25) => PC_BUS_25_port, 
                           PC_BUS(24) => PC_BUS_24_port, PC_BUS(23) => 
                           PC_BUS_23_port, PC_BUS(22) => PC_BUS_22_port, 
                           PC_BUS(21) => PC_BUS_21_port, PC_BUS(20) => 
                           PC_BUS_20_port, PC_BUS(19) => PC_BUS_19_port, 
                           PC_BUS(18) => PC_BUS_18_port, PC_BUS(17) => 
                           PC_BUS_17_port, PC_BUS(16) => PC_BUS_16_port, 
                           PC_BUS(15) => PC_BUS_15_port, PC_BUS(14) => 
                           PC_BUS_14_port, PC_BUS(13) => PC_BUS_13_port, 
                           PC_BUS(12) => PC_BUS_12_port, PC_BUS(11) => 
                           PC_BUS_11_port, PC_BUS(10) => PC_BUS_10_port, 
                           PC_BUS(9) => PC_BUS_9_port, PC_BUS(8) => 
                           PC_BUS_8_port, PC_BUS(7) => PC_BUS_7_port, PC_BUS(6)
                           => PC_BUS_6_port, PC_BUS(5) => PC_BUS_5_port, 
                           PC_BUS(4) => PC_BUS_4_port, PC_BUS(3) => 
                           PC_BUS_3_port, PC_BUS(2) => PC_BUS_2_port, PC_BUS(1)
                           => PC_BUS_1_port, PC_BUS(0) => PC_BUS_0_port);
   CU : dlx_cu port map( Clk => CLK, Rst => RST, IR_IN(31) => I_DATA(31), 
                           IR_IN(30) => I_DATA(30), IR_IN(29) => I_DATA(29), 
                           IR_IN(28) => I_DATA(28), IR_IN(27) => I_DATA(27), 
                           IR_IN(26) => I_DATA(26), IR_IN(25) => I_DATA(25), 
                           IR_IN(24) => I_DATA(24), IR_IN(23) => I_DATA(23), 
                           IR_IN(22) => I_DATA(22), IR_IN(21) => I_DATA(21), 
                           IR_IN(20) => I_DATA(20), IR_IN(19) => I_DATA(19), 
                           IR_IN(18) => I_DATA(18), IR_IN(17) => I_DATA(17), 
                           IR_IN(16) => I_DATA(16), IR_IN(15) => I_DATA(15), 
                           IR_IN(14) => I_DATA(14), IR_IN(13) => I_DATA(13), 
                           IR_IN(12) => I_DATA(12), IR_IN(11) => I_DATA(11), 
                           IR_IN(10) => I_DATA(10), IR_IN(9) => I_DATA(9), 
                           IR_IN(8) => I_DATA(8), IR_IN(7) => I_DATA(7), 
                           IR_IN(6) => I_DATA(6), IR_IN(5) => I_DATA(5), 
                           IR_IN(4) => I_DATA(4), IR_IN(3) => I_DATA(3), 
                           IR_IN(2) => I_DATA(2), IR_IN(1) => I_DATA(1), 
                           IR_IN(0) => I_DATA(0), IR_LATCH_EN => n_2424, 
                           NPC_LATCH_EN => n_2425, RegA_LATCH_EN => n_2426, 
                           RegB_LATCH_EN => n_2427, RegIMM_LATCH_EN => n_2428, 
                           SIGNED_IMM => n_2429, MUXA_SEL => n_2430, MUXB_SEL 
                           => n_2431, ALU_OUTREG_EN => n_2432, EQ_COND => 
                           n_2433, IS_JUMP => n_2434, ALU_OPCODE(0) => 
                           ALU_OPCODE_3_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_2_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_1_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_0_port, DRAM_WE => n_2435, LMD_LATCH_EN 
                           => n_2436, JUMP_EN => n_2437, PC_LATCH_EN => n_2438,
                           IS_JAL => n_2439, WB_MUX_SEL => n_2440, RF_WE => 
                           n_2441);

end SYN_DLX_RTL;
