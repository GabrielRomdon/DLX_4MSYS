
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOpType is (NOP, ADDS, SUBS, ANDS, ORS, XORS, SLE, SGE, SNE, SRLS, SLLS)
   ;
attribute ENUM_ENCODING of aluOpType : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOpType(arg : in std_logic_vector( 1 to 4 )) 
               return aluOpType;
   function aluOpType_to_std_logic_vector(arg : in aluOpType) return 
               std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOpType(arg : in std_logic_vector( 1 to 4 )) 
   return aluOpType is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "0000" => return NOP;
         when "0001" => return ADDS;
         when "0010" => return SUBS;
         when "0011" => return ANDS;
         when "0100" => return ORS;
         when "0101" => return XORS;
         when "0110" => return SLE;
         when "0111" => return SGE;
         when "1000" => return SNE;
         when "1001" => return SRLS;
         when "1010" => return SLLS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOpType_to_std_logic_vector(arg : in aluOpType) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "0000";
         when ADDS => return "0001";
         when SUBS => return "0010";
         when ANDS => return "0011";
         when ORS => return "0100";
         when XORS => return "0101";
         when SLE => return "0110";
         when SGE => return "0111";
         when SNE => return "1000";
         when SRLS => return "1001";
         when SLLS => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_N32_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end ADDER_N32_DW01_add_0;

architecture SYN_rpl of ADDER_N32_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, SUM_3_port,
      SUM_4_port, SUM_5_port, SUM_6_port, SUM_7_port, SUM_8_port, SUM_9_port, 
      SUM_10_port, SUM_11_port, SUM_12_port, SUM_13_port, SUM_14_port, 
      SUM_15_port, SUM_16_port, SUM_17_port, SUM_18_port, SUM_19_port, 
      SUM_20_port, SUM_21_port, SUM_22_port, SUM_23_port, SUM_24_port, 
      SUM_25_port, SUM_26_port, SUM_27_port, SUM_28_port, SUM_29_port, 
      SUM_30_port, SUM_31_port, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : AND2_X1 port map( A1 => A(9), A2 => n7, ZN => n1);
   U2 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n2);
   U3 : AND2_X1 port map( A1 => A(4), A2 => n2, ZN => n3);
   U4 : AND2_X1 port map( A1 => A(5), A2 => n3, ZN => n4);
   U5 : AND2_X1 port map( A1 => A(6), A2 => n4, ZN => n5);
   U6 : AND2_X1 port map( A1 => A(7), A2 => n5, ZN => n6);
   U7 : AND2_X1 port map( A1 => A(8), A2 => n6, ZN => n7);
   U8 : AND2_X1 port map( A1 => A(10), A2 => n1, ZN => n8);
   U9 : AND2_X1 port map( A1 => A(11), A2 => n8, ZN => n9);
   U10 : AND2_X1 port map( A1 => A(12), A2 => n9, ZN => n10);
   U11 : AND2_X1 port map( A1 => A(13), A2 => n10, ZN => n11);
   U12 : AND2_X1 port map( A1 => A(14), A2 => n11, ZN => n12);
   U13 : AND2_X1 port map( A1 => A(15), A2 => n12, ZN => n13);
   U14 : AND2_X1 port map( A1 => A(16), A2 => n13, ZN => n14);
   U15 : AND2_X1 port map( A1 => A(17), A2 => n14, ZN => n15);
   U16 : AND2_X1 port map( A1 => A(18), A2 => n15, ZN => n16);
   U17 : AND2_X1 port map( A1 => A(19), A2 => n16, ZN => n17);
   U18 : AND2_X1 port map( A1 => A(20), A2 => n17, ZN => n18);
   U19 : AND2_X1 port map( A1 => A(21), A2 => n18, ZN => n19);
   U20 : AND2_X1 port map( A1 => A(22), A2 => n19, ZN => n20);
   U21 : AND2_X1 port map( A1 => A(23), A2 => n20, ZN => n21);
   U22 : AND2_X1 port map( A1 => A(24), A2 => n21, ZN => n22);
   U23 : AND2_X1 port map( A1 => A(25), A2 => n22, ZN => n23);
   U24 : AND2_X1 port map( A1 => A(26), A2 => n23, ZN => n24);
   U25 : AND2_X1 port map( A1 => A(27), A2 => n24, ZN => n25);
   U26 : AND2_X1 port map( A1 => A(28), A2 => n25, ZN => n26);
   U27 : AND2_X1 port map( A1 => A(29), A2 => n26, ZN => n27);
   U28 : AND2_X1 port map( A1 => A(30), A2 => n27, ZN => n28);
   U29 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U30 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U31 : XOR2_X1 port map( A => A(4), B => n2, Z => SUM_4_port);
   U32 : XOR2_X1 port map( A => A(5), B => n3, Z => SUM_5_port);
   U33 : XOR2_X1 port map( A => A(6), B => n4, Z => SUM_6_port);
   U34 : XOR2_X1 port map( A => A(7), B => n5, Z => SUM_7_port);
   U35 : XOR2_X1 port map( A => A(8), B => n6, Z => SUM_8_port);
   U36 : XOR2_X1 port map( A => A(9), B => n7, Z => SUM_9_port);
   U37 : XOR2_X1 port map( A => A(10), B => n1, Z => SUM_10_port);
   U38 : XOR2_X1 port map( A => A(11), B => n8, Z => SUM_11_port);
   U39 : XOR2_X1 port map( A => A(12), B => n9, Z => SUM_12_port);
   U40 : XOR2_X1 port map( A => A(13), B => n10, Z => SUM_13_port);
   U41 : XOR2_X1 port map( A => A(14), B => n11, Z => SUM_14_port);
   U42 : XOR2_X1 port map( A => A(15), B => n12, Z => SUM_15_port);
   U43 : XOR2_X1 port map( A => A(16), B => n13, Z => SUM_16_port);
   U44 : XOR2_X1 port map( A => A(17), B => n14, Z => SUM_17_port);
   U45 : XOR2_X1 port map( A => A(18), B => n15, Z => SUM_18_port);
   U46 : XOR2_X1 port map( A => A(19), B => n16, Z => SUM_19_port);
   U47 : XOR2_X1 port map( A => A(20), B => n17, Z => SUM_20_port);
   U48 : XOR2_X1 port map( A => A(21), B => n18, Z => SUM_21_port);
   U49 : XOR2_X1 port map( A => A(22), B => n19, Z => SUM_22_port);
   U50 : XOR2_X1 port map( A => A(23), B => n20, Z => SUM_23_port);
   U51 : XOR2_X1 port map( A => A(24), B => n21, Z => SUM_24_port);
   U52 : XOR2_X1 port map( A => A(25), B => n22, Z => SUM_25_port);
   U53 : XOR2_X1 port map( A => A(26), B => n23, Z => SUM_26_port);
   U54 : XOR2_X1 port map( A => A(27), B => n24, Z => SUM_27_port);
   U55 : XOR2_X1 port map( A => A(28), B => n25, Z => SUM_28_port);
   U56 : XOR2_X1 port map( A => A(29), B => n26, Z => SUM_29_port);
   U57 : XOR2_X1 port map( A => A(30), B => n27, Z => SUM_30_port);
   U58 : XOR2_X1 port map( A => A(31), B => n28, Z => SUM_31_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end ALU_N32_DW01_cmp6_0;

architecture SYN_rpl of ALU_N32_DW01_cmp6_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal GE_port, LE_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208 : 
      std_logic;

begin
   LE <= LE_port;
   GE <= GE_port;
   
   U1 : INV_X1 port map( A => n135, ZN => n27);
   U2 : INV_X1 port map( A => n125, ZN => n23);
   U3 : INV_X1 port map( A => n115, ZN => n19);
   U4 : INV_X1 port map( A => n85, ZN => n7);
   U5 : INV_X1 port map( A => n105, ZN => n15);
   U6 : INV_X1 port map( A => n95, ZN => n11);
   U7 : INV_X1 port map( A => n131, ZN => n28);
   U8 : INV_X1 port map( A => n121, ZN => n24);
   U9 : INV_X1 port map( A => n111, ZN => n20);
   U10 : INV_X1 port map( A => n101, ZN => n16);
   U11 : INV_X1 port map( A => n91, ZN => n12);
   U12 : INV_X1 port map( A => n81, ZN => n8);
   U13 : INV_X1 port map( A => n140, ZN => n31);
   U14 : INV_X1 port map( A => n114, ZN => n21);
   U15 : INV_X1 port map( A => n130, ZN => n26);
   U16 : INV_X1 port map( A => n100, ZN => n14);
   U17 : INV_X1 port map( A => n84, ZN => n9);
   U18 : INV_X1 port map( A => n134, ZN => n29);
   U19 : INV_X1 port map( A => n104, ZN => n17);
   U20 : INV_X1 port map( A => n120, ZN => n22);
   U21 : INV_X1 port map( A => n90, ZN => n10);
   U22 : INV_X1 port map( A => n75, ZN => n5);
   U23 : INV_X1 port map( A => n139, ZN => n30);
   U24 : INV_X1 port map( A => n110, ZN => n18);
   U25 : INV_X1 port map( A => n80, ZN => n6);
   U26 : INV_X1 port map( A => n124, ZN => n25);
   U27 : INV_X1 port map( A => n94, ZN => n13);
   U28 : INV_X1 port map( A => B(2), ZN => n63);
   U29 : INV_X1 port map( A => B(0), ZN => n64);
   U30 : INV_X1 port map( A => n206, ZN => n32);
   U31 : INV_X1 port map( A => n65, ZN => LE_port);
   U32 : INV_X1 port map( A => A(31), ZN => n3);
   U33 : INV_X1 port map( A => A(1), ZN => n33);
   U34 : INV_X1 port map( A => n144, ZN => n34);
   U35 : INV_X1 port map( A => B(3), ZN => n62);
   U36 : INV_X1 port map( A => A(30), ZN => n4);
   U37 : INV_X1 port map( A => B(4), ZN => n61);
   U38 : INV_X1 port map( A => B(6), ZN => n59);
   U39 : INV_X1 port map( A => B(10), ZN => n55);
   U40 : INV_X1 port map( A => B(14), ZN => n51);
   U41 : INV_X1 port map( A => B(18), ZN => n47);
   U42 : INV_X1 port map( A => B(22), ZN => n43);
   U43 : INV_X1 port map( A => B(26), ZN => n39);
   U44 : INV_X1 port map( A => B(30), ZN => n35);
   U45 : INV_X1 port map( A => B(8), ZN => n57);
   U46 : INV_X1 port map( A => B(12), ZN => n53);
   U47 : INV_X1 port map( A => B(5), ZN => n60);
   U48 : INV_X1 port map( A => B(16), ZN => n49);
   U49 : INV_X1 port map( A => B(9), ZN => n56);
   U50 : INV_X1 port map( A => B(13), ZN => n52);
   U51 : INV_X1 port map( A => B(20), ZN => n45);
   U52 : INV_X1 port map( A => B(17), ZN => n48);
   U53 : INV_X1 port map( A => B(21), ZN => n44);
   U54 : INV_X1 port map( A => B(24), ZN => n41);
   U55 : INV_X1 port map( A => B(25), ZN => n40);
   U56 : INV_X1 port map( A => B(28), ZN => n37);
   U57 : INV_X1 port map( A => B(29), ZN => n36);
   U58 : INV_X1 port map( A => B(7), ZN => n58);
   U59 : INV_X1 port map( A => B(11), ZN => n54);
   U60 : INV_X1 port map( A => B(15), ZN => n50);
   U61 : INV_X1 port map( A => B(19), ZN => n46);
   U62 : INV_X1 port map( A => B(23), ZN => n42);
   U63 : INV_X1 port map( A => B(27), ZN => n38);
   U64 : INV_X1 port map( A => n159, ZN => GE_port);
   U65 : NAND2_X1 port map( A1 => GE_port, A2 => LE_port, ZN => NE);
   U66 : OAI21_X1 port map( B1 => n66, B2 => n67, A => n68, ZN => n65);
   U67 : MUX2_X1 port map( A => n69, B => n70, S => n3, Z => n68);
   U68 : NAND2_X1 port map( A1 => TC, A2 => B(31), ZN => n70);
   U69 : OR2_X1 port map( A1 => B(31), A2 => TC, ZN => n69);
   U70 : AOI22_X1 port map( A1 => A(30), A2 => n35, B1 => n71, B2 => n72, ZN =>
                           n66);
   U71 : AOI21_X1 port map( B1 => n73, B2 => n74, A => n75, ZN => n71);
   U72 : OAI211_X1 port map( C1 => n76, C2 => n77, A => n78, B => n79, ZN => 
                           n74);
   U73 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => n77);
   U74 : AOI211_X1 port map( C1 => n82, C2 => n83, A => n7, B => n84, ZN => n76
                           );
   U75 : OAI211_X1 port map( C1 => n86, C2 => n87, A => n88, B => n89, ZN => 
                           n83);
   U76 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => n87);
   U77 : AOI211_X1 port map( C1 => n92, C2 => n93, A => n11, B => n94, ZN => 
                           n86);
   U78 : OAI211_X1 port map( C1 => n96, C2 => n97, A => n98, B => n99, ZN => 
                           n93);
   U79 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => n97);
   U80 : AOI211_X1 port map( C1 => n102, C2 => n103, A => n15, B => n104, ZN =>
                           n96);
   U81 : OAI211_X1 port map( C1 => n106, C2 => n107, A => n108, B => n109, ZN 
                           => n103);
   U82 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => n107);
   U83 : AOI211_X1 port map( C1 => n112, C2 => n113, A => n19, B => n114, ZN =>
                           n106);
   U84 : OAI211_X1 port map( C1 => n116, C2 => n117, A => n118, B => n119, ZN 
                           => n113);
   U85 : NAND2_X1 port map( A1 => n120, A2 => n121, ZN => n117);
   U86 : AOI211_X1 port map( C1 => n122, C2 => n123, A => n23, B => n124, ZN =>
                           n116);
   U87 : OAI211_X1 port map( C1 => n126, C2 => n127, A => n128, B => n129, ZN 
                           => n123);
   U88 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => n127);
   U89 : AOI211_X1 port map( C1 => n132, C2 => n133, A => n27, B => n134, ZN =>
                           n126);
   U90 : NAND3_X1 port map( A1 => n136, A2 => n137, A3 => n138, ZN => n133);
   U91 : NAND3_X1 port map( A1 => n139, A2 => n140, A3 => n141, ZN => n136);
   U92 : OAI211_X1 port map( C1 => A(1), C2 => n34, A => n142, B => n143, ZN =>
                           n141);
   U93 : OAI21_X1 port map( B1 => n33, B2 => n144, A => B(1), ZN => n142);
   U94 : NAND2_X1 port map( A1 => A(0), A2 => n64, ZN => n144);
   U95 : NOR2_X1 port map( A1 => n145, A2 => n146, ZN => n132);
   U96 : NOR2_X1 port map( A1 => n147, A2 => n148, ZN => n122);
   U97 : NOR2_X1 port map( A1 => n149, A2 => n150, ZN => n112);
   U98 : NOR2_X1 port map( A1 => n151, A2 => n152, ZN => n102);
   U99 : NOR2_X1 port map( A1 => n153, A2 => n154, ZN => n92);
   U100 : NOR2_X1 port map( A1 => n155, A2 => n156, ZN => n82);
   U101 : NOR2_X1 port map( A1 => n157, A2 => n158, ZN => n73);
   U102 : OAI21_X1 port map( B1 => n160, B2 => n67, A => n161, ZN => n159);
   U103 : MUX2_X1 port map( A => n162, B => n163, S => TC, Z => n161);
   U104 : OR2_X1 port map( A1 => n3, A2 => B(31), ZN => n163);
   U105 : NAND2_X1 port map( A1 => B(31), A2 => n3, ZN => n162);
   U106 : XNOR2_X1 port map( A => n3, B => B(31), ZN => n67);
   U107 : AOI22_X1 port map( A1 => B(30), A2 => n4, B1 => n164, B2 => n72, ZN 
                           => n160);
   U108 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n72);
   U109 : AOI21_X1 port map( B1 => n165, B2 => n5, A => n158, ZN => n164);
   U110 : AND2_X1 port map( A1 => A(29), A2 => n36, ZN => n158);
   U111 : NOR2_X1 port map( A1 => n36, A2 => A(29), ZN => n75);
   U112 : AOI21_X1 port map( B1 => n166, B2 => n79, A => n167, ZN => n165);
   U113 : NOR2_X1 port map( A1 => n167, A2 => n157, ZN => n79);
   U114 : AND2_X1 port map( A1 => A(28), A2 => n37, ZN => n157);
   U115 : NOR2_X1 port map( A1 => n37, A2 => A(28), ZN => n167);
   U116 : AOI21_X1 port map( B1 => n168, B2 => n78, A => n6, ZN => n166);
   U117 : NAND2_X1 port map( A1 => A(27), A2 => n38, ZN => n80);
   U118 : OR2_X1 port map( A1 => n38, A2 => A(27), ZN => n78);
   U119 : AOI21_X1 port map( B1 => n169, B2 => n85, A => n170, ZN => n168);
   U120 : NOR2_X1 port map( A1 => n170, A2 => n8, ZN => n85);
   U121 : NAND2_X1 port map( A1 => A(26), A2 => n39, ZN => n81);
   U122 : NOR2_X1 port map( A1 => n39, A2 => A(26), ZN => n170);
   U123 : AOI21_X1 port map( B1 => n171, B2 => n9, A => n156, ZN => n169);
   U124 : AND2_X1 port map( A1 => A(25), A2 => n40, ZN => n156);
   U125 : NOR2_X1 port map( A1 => n40, A2 => A(25), ZN => n84);
   U126 : AOI21_X1 port map( B1 => n172, B2 => n89, A => n173, ZN => n171);
   U127 : NOR2_X1 port map( A1 => n173, A2 => n155, ZN => n89);
   U128 : AND2_X1 port map( A1 => A(24), A2 => n41, ZN => n155);
   U129 : NOR2_X1 port map( A1 => n41, A2 => A(24), ZN => n173);
   U130 : AOI21_X1 port map( B1 => n174, B2 => n88, A => n10, ZN => n172);
   U131 : NAND2_X1 port map( A1 => A(23), A2 => n42, ZN => n90);
   U132 : OR2_X1 port map( A1 => n42, A2 => A(23), ZN => n88);
   U133 : AOI21_X1 port map( B1 => n175, B2 => n95, A => n176, ZN => n174);
   U134 : NOR2_X1 port map( A1 => n176, A2 => n12, ZN => n95);
   U135 : NAND2_X1 port map( A1 => A(22), A2 => n43, ZN => n91);
   U136 : NOR2_X1 port map( A1 => n43, A2 => A(22), ZN => n176);
   U137 : AOI21_X1 port map( B1 => n177, B2 => n13, A => n154, ZN => n175);
   U138 : AND2_X1 port map( A1 => A(21), A2 => n44, ZN => n154);
   U139 : NOR2_X1 port map( A1 => n44, A2 => A(21), ZN => n94);
   U140 : AOI21_X1 port map( B1 => n178, B2 => n99, A => n179, ZN => n177);
   U141 : NOR2_X1 port map( A1 => n179, A2 => n153, ZN => n99);
   U142 : AND2_X1 port map( A1 => A(20), A2 => n45, ZN => n153);
   U143 : NOR2_X1 port map( A1 => n45, A2 => A(20), ZN => n179);
   U144 : AOI21_X1 port map( B1 => n180, B2 => n98, A => n14, ZN => n178);
   U145 : NAND2_X1 port map( A1 => A(19), A2 => n46, ZN => n100);
   U146 : OR2_X1 port map( A1 => n46, A2 => A(19), ZN => n98);
   U147 : AOI21_X1 port map( B1 => n181, B2 => n105, A => n182, ZN => n180);
   U148 : NOR2_X1 port map( A1 => n182, A2 => n16, ZN => n105);
   U149 : NAND2_X1 port map( A1 => A(18), A2 => n47, ZN => n101);
   U150 : NOR2_X1 port map( A1 => n47, A2 => A(18), ZN => n182);
   U151 : AOI21_X1 port map( B1 => n183, B2 => n17, A => n152, ZN => n181);
   U152 : AND2_X1 port map( A1 => A(17), A2 => n48, ZN => n152);
   U153 : NOR2_X1 port map( A1 => n48, A2 => A(17), ZN => n104);
   U154 : AOI21_X1 port map( B1 => n184, B2 => n109, A => n185, ZN => n183);
   U155 : NOR2_X1 port map( A1 => n185, A2 => n151, ZN => n109);
   U156 : AND2_X1 port map( A1 => A(16), A2 => n49, ZN => n151);
   U157 : NOR2_X1 port map( A1 => n49, A2 => A(16), ZN => n185);
   U158 : AOI21_X1 port map( B1 => n186, B2 => n108, A => n18, ZN => n184);
   U159 : NAND2_X1 port map( A1 => A(15), A2 => n50, ZN => n110);
   U160 : OR2_X1 port map( A1 => n50, A2 => A(15), ZN => n108);
   U161 : AOI21_X1 port map( B1 => n187, B2 => n115, A => n188, ZN => n186);
   U162 : NOR2_X1 port map( A1 => n188, A2 => n20, ZN => n115);
   U163 : NAND2_X1 port map( A1 => A(14), A2 => n51, ZN => n111);
   U164 : NOR2_X1 port map( A1 => n51, A2 => A(14), ZN => n188);
   U165 : AOI21_X1 port map( B1 => n189, B2 => n21, A => n150, ZN => n187);
   U166 : AND2_X1 port map( A1 => A(13), A2 => n52, ZN => n150);
   U167 : NOR2_X1 port map( A1 => n52, A2 => A(13), ZN => n114);
   U168 : AOI21_X1 port map( B1 => n190, B2 => n119, A => n191, ZN => n189);
   U169 : NOR2_X1 port map( A1 => n191, A2 => n149, ZN => n119);
   U170 : AND2_X1 port map( A1 => A(12), A2 => n53, ZN => n149);
   U171 : NOR2_X1 port map( A1 => n53, A2 => A(12), ZN => n191);
   U172 : AOI21_X1 port map( B1 => n192, B2 => n118, A => n22, ZN => n190);
   U173 : NAND2_X1 port map( A1 => A(11), A2 => n54, ZN => n120);
   U174 : OR2_X1 port map( A1 => n54, A2 => A(11), ZN => n118);
   U175 : AOI21_X1 port map( B1 => n193, B2 => n125, A => n194, ZN => n192);
   U176 : NOR2_X1 port map( A1 => n194, A2 => n24, ZN => n125);
   U177 : NAND2_X1 port map( A1 => A(10), A2 => n55, ZN => n121);
   U178 : NOR2_X1 port map( A1 => n55, A2 => A(10), ZN => n194);
   U179 : AOI21_X1 port map( B1 => n195, B2 => n25, A => n148, ZN => n193);
   U180 : AND2_X1 port map( A1 => A(9), A2 => n56, ZN => n148);
   U181 : NOR2_X1 port map( A1 => n56, A2 => A(9), ZN => n124);
   U182 : AOI21_X1 port map( B1 => n196, B2 => n129, A => n197, ZN => n195);
   U183 : NOR2_X1 port map( A1 => n197, A2 => n147, ZN => n129);
   U184 : AND2_X1 port map( A1 => A(8), A2 => n57, ZN => n147);
   U185 : NOR2_X1 port map( A1 => n57, A2 => A(8), ZN => n197);
   U186 : AOI21_X1 port map( B1 => n198, B2 => n128, A => n26, ZN => n196);
   U187 : NAND2_X1 port map( A1 => A(7), A2 => n58, ZN => n130);
   U188 : OR2_X1 port map( A1 => n58, A2 => A(7), ZN => n128);
   U189 : AOI21_X1 port map( B1 => n199, B2 => n135, A => n200, ZN => n198);
   U190 : NOR2_X1 port map( A1 => n200, A2 => n28, ZN => n135);
   U191 : NAND2_X1 port map( A1 => A(6), A2 => n59, ZN => n131);
   U192 : NOR2_X1 port map( A1 => n59, A2 => A(6), ZN => n200);
   U193 : AOI21_X1 port map( B1 => n201, B2 => n29, A => n146, ZN => n199);
   U194 : AND2_X1 port map( A1 => A(5), A2 => n60, ZN => n146);
   U195 : NOR2_X1 port map( A1 => n60, A2 => A(5), ZN => n134);
   U196 : AOI21_X1 port map( B1 => n202, B2 => n138, A => n203, ZN => n201);
   U197 : NOR2_X1 port map( A1 => n203, A2 => n145, ZN => n138);
   U198 : AND2_X1 port map( A1 => A(4), A2 => n61, ZN => n145);
   U199 : NOR2_X1 port map( A1 => n61, A2 => A(4), ZN => n203);
   U200 : AOI21_X1 port map( B1 => n204, B2 => n137, A => n30, ZN => n202);
   U201 : NAND2_X1 port map( A1 => A(3), A2 => n62, ZN => n139);
   U202 : OR2_X1 port map( A1 => n62, A2 => A(3), ZN => n137);
   U203 : AOI21_X1 port map( B1 => n32, B2 => n143, A => n205, ZN => n204);
   U204 : NOR2_X1 port map( A1 => n205, A2 => n31, ZN => n143);
   U205 : NAND2_X1 port map( A1 => A(2), A2 => n63, ZN => n140);
   U206 : NOR2_X1 port map( A1 => n63, A2 => A(2), ZN => n205);
   U207 : OAI22_X1 port map( A1 => n207, A2 => B(1), B1 => n33, B2 => n208, ZN 
                           => n206);
   U208 : AND2_X1 port map( A1 => n208, A2 => n33, ZN => n207);
   U209 : NOR2_X1 port map( A1 => n64, A2 => A(0), ZN => n208);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_addsub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in std_logic;
         SUM : out std_logic_vector (31 downto 0);  CO : out std_logic);

end ALU_N32_DW01_addsub_0;

architecture SYN_rpl of ALU_N32_DW01_addsub_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, B_AS_31_port, 
      B_AS_30_port, B_AS_29_port, B_AS_28_port, B_AS_27_port, B_AS_26_port, 
      B_AS_25_port, B_AS_24_port, B_AS_23_port, B_AS_22_port, B_AS_21_port, 
      B_AS_20_port, B_AS_19_port, B_AS_18_port, B_AS_17_port, B_AS_16_port, 
      B_AS_15_port, B_AS_14_port, B_AS_13_port, B_AS_12_port, B_AS_11_port, 
      B_AS_10_port, B_AS_9_port, B_AS_8_port, B_AS_7_port, B_AS_6_port, 
      B_AS_5_port, B_AS_4_port, B_AS_3_port, B_AS_2_port, B_AS_1_port, 
      B_AS_0_port, n_1039 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B_AS_31_port, CI => carry_31_port, 
                           CO => n_1039, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B_AS_30_port, CI => carry_30_port, 
                           CO => carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B_AS_29_port, CI => carry_29_port, 
                           CO => carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B_AS_28_port, CI => carry_28_port, 
                           CO => carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B_AS_27_port, CI => carry_27_port, 
                           CO => carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B_AS_26_port, CI => carry_26_port, 
                           CO => carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B_AS_25_port, CI => carry_25_port, 
                           CO => carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B_AS_24_port, CI => carry_24_port, 
                           CO => carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B_AS_23_port, CI => carry_23_port, 
                           CO => carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B_AS_22_port, CI => carry_22_port, 
                           CO => carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B_AS_21_port, CI => carry_21_port, 
                           CO => carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B_AS_20_port, CI => carry_20_port, 
                           CO => carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B_AS_19_port, CI => carry_19_port, 
                           CO => carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B_AS_18_port, CI => carry_18_port, 
                           CO => carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B_AS_17_port, CI => carry_17_port, 
                           CO => carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B_AS_16_port, CI => carry_16_port, 
                           CO => carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B_AS_15_port, CI => carry_15_port, 
                           CO => carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B_AS_14_port, CI => carry_14_port, 
                           CO => carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B_AS_13_port, CI => carry_13_port, 
                           CO => carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B_AS_12_port, CI => carry_12_port, 
                           CO => carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B_AS_11_port, CI => carry_11_port, 
                           CO => carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B_AS_10_port, CI => carry_10_port, 
                           CO => carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B_AS_9_port, CI => carry_9_port, CO 
                           => carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B_AS_8_port, CI => carry_8_port, CO 
                           => carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B_AS_7_port, CI => carry_7_port, CO 
                           => carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B_AS_6_port, CI => carry_6_port, CO 
                           => carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B_AS_5_port, CI => carry_5_port, CO 
                           => carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B_AS_4_port, CI => carry_4_port, CO 
                           => carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B_AS_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B_AS_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B_AS_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_AS_9_port);
   U2 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_AS_8_port);
   U3 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_AS_7_port);
   U4 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_AS_6_port);
   U5 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_AS_5_port);
   U6 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_AS_4_port);
   U7 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_AS_3_port);
   U8 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_AS_31_port);
   U9 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_AS_30_port);
   U10 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_AS_2_port);
   U11 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_AS_29_port);
   U12 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_AS_28_port);
   U13 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_AS_27_port);
   U14 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_AS_26_port);
   U15 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_AS_25_port);
   U16 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_AS_24_port);
   U17 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_AS_23_port);
   U18 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_AS_22_port);
   U19 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_AS_21_port);
   U20 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_AS_20_port);
   U21 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_AS_1_port);
   U22 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_AS_19_port);
   U23 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_AS_18_port);
   U24 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_AS_17_port);
   U25 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_AS_16_port);
   U26 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_AS_15_port);
   U27 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_AS_14_port);
   U28 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_AS_13_port);
   U29 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_AS_12_port);
   U30 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_AS_11_port);
   U31 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_AS_10_port);
   U32 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_31 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_31;

architecture SYN_BEHAVIOUR of NAND4_31 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_30 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_30;

architecture SYN_BEHAVIOUR of NAND4_30 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_29 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_29;

architecture SYN_BEHAVIOUR of NAND4_29 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_28 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_28;

architecture SYN_BEHAVIOUR of NAND4_28 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_27 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_27;

architecture SYN_BEHAVIOUR of NAND4_27 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_26 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_26;

architecture SYN_BEHAVIOUR of NAND4_26 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_25 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_25;

architecture SYN_BEHAVIOUR of NAND4_25 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_24 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_24;

architecture SYN_BEHAVIOUR of NAND4_24 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_23 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_23;

architecture SYN_BEHAVIOUR of NAND4_23 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_22 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_22;

architecture SYN_BEHAVIOUR of NAND4_22 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_21 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_21;

architecture SYN_BEHAVIOUR of NAND4_21 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_20 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_20;

architecture SYN_BEHAVIOUR of NAND4_20 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_19 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_19;

architecture SYN_BEHAVIOUR of NAND4_19 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_18 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_18;

architecture SYN_BEHAVIOUR of NAND4_18 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_17 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_17;

architecture SYN_BEHAVIOUR of NAND4_17 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_16 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_16;

architecture SYN_BEHAVIOUR of NAND4_16 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_15 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_15;

architecture SYN_BEHAVIOUR of NAND4_15 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_14 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_14;

architecture SYN_BEHAVIOUR of NAND4_14 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_13 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_13;

architecture SYN_BEHAVIOUR of NAND4_13 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_12 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_12;

architecture SYN_BEHAVIOUR of NAND4_12 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_11 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_11;

architecture SYN_BEHAVIOUR of NAND4_11 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_10 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_10;

architecture SYN_BEHAVIOUR of NAND4_10 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_9 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_9;

architecture SYN_BEHAVIOUR of NAND4_9 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_8 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_8;

architecture SYN_BEHAVIOUR of NAND4_8 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_7 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_7;

architecture SYN_BEHAVIOUR of NAND4_7 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_6 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_6;

architecture SYN_BEHAVIOUR of NAND4_6 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_5 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_5;

architecture SYN_BEHAVIOUR of NAND4_5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_4 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_4;

architecture SYN_BEHAVIOUR of NAND4_4 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_3 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_3;

architecture SYN_BEHAVIOUR of NAND4_3 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_2 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_2;

architecture SYN_BEHAVIOUR of NAND4_2 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_1 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_1;

architecture SYN_BEHAVIOUR of NAND4_1 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_127 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_127;

architecture SYN_BEHAVIOUR of NAND3_127 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_126 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_126;

architecture SYN_BEHAVIOUR of NAND3_126 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_125 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_125;

architecture SYN_BEHAVIOUR of NAND3_125 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_124 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_124;

architecture SYN_BEHAVIOUR of NAND3_124 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_123 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_123;

architecture SYN_BEHAVIOUR of NAND3_123 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_122 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_122;

architecture SYN_BEHAVIOUR of NAND3_122 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_121 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_121;

architecture SYN_BEHAVIOUR of NAND3_121 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_120 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_120;

architecture SYN_BEHAVIOUR of NAND3_120 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_119 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_119;

architecture SYN_BEHAVIOUR of NAND3_119 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_118 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_118;

architecture SYN_BEHAVIOUR of NAND3_118 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_117 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_117;

architecture SYN_BEHAVIOUR of NAND3_117 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_116 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_116;

architecture SYN_BEHAVIOUR of NAND3_116 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_115 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_115;

architecture SYN_BEHAVIOUR of NAND3_115 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_114 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_114;

architecture SYN_BEHAVIOUR of NAND3_114 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_113 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_113;

architecture SYN_BEHAVIOUR of NAND3_113 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_112 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_112;

architecture SYN_BEHAVIOUR of NAND3_112 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_111 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_111;

architecture SYN_BEHAVIOUR of NAND3_111 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_110 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_110;

architecture SYN_BEHAVIOUR of NAND3_110 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_109 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_109;

architecture SYN_BEHAVIOUR of NAND3_109 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_108 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_108;

architecture SYN_BEHAVIOUR of NAND3_108 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_107 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_107;

architecture SYN_BEHAVIOUR of NAND3_107 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_106 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_106;

architecture SYN_BEHAVIOUR of NAND3_106 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_105 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_105;

architecture SYN_BEHAVIOUR of NAND3_105 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_104 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_104;

architecture SYN_BEHAVIOUR of NAND3_104 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_103 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_103;

architecture SYN_BEHAVIOUR of NAND3_103 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_102 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_102;

architecture SYN_BEHAVIOUR of NAND3_102 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_101 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_101;

architecture SYN_BEHAVIOUR of NAND3_101 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_100 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_100;

architecture SYN_BEHAVIOUR of NAND3_100 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_99 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_99;

architecture SYN_BEHAVIOUR of NAND3_99 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_98 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_98;

architecture SYN_BEHAVIOUR of NAND3_98 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_97 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_97;

architecture SYN_BEHAVIOUR of NAND3_97 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_96 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_96;

architecture SYN_BEHAVIOUR of NAND3_96 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_95 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_95;

architecture SYN_BEHAVIOUR of NAND3_95 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_94 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_94;

architecture SYN_BEHAVIOUR of NAND3_94 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_93 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_93;

architecture SYN_BEHAVIOUR of NAND3_93 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_92 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_92;

architecture SYN_BEHAVIOUR of NAND3_92 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_91 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_91;

architecture SYN_BEHAVIOUR of NAND3_91 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_90 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_90;

architecture SYN_BEHAVIOUR of NAND3_90 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_89 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_89;

architecture SYN_BEHAVIOUR of NAND3_89 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_88 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_88;

architecture SYN_BEHAVIOUR of NAND3_88 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_87 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_87;

architecture SYN_BEHAVIOUR of NAND3_87 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_86 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_86;

architecture SYN_BEHAVIOUR of NAND3_86 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_85 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_85;

architecture SYN_BEHAVIOUR of NAND3_85 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_84 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_84;

architecture SYN_BEHAVIOUR of NAND3_84 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_83 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_83;

architecture SYN_BEHAVIOUR of NAND3_83 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_82 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_82;

architecture SYN_BEHAVIOUR of NAND3_82 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_81 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_81;

architecture SYN_BEHAVIOUR of NAND3_81 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_80 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_80;

architecture SYN_BEHAVIOUR of NAND3_80 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_79 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_79;

architecture SYN_BEHAVIOUR of NAND3_79 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_78 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_78;

architecture SYN_BEHAVIOUR of NAND3_78 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_77 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_77;

architecture SYN_BEHAVIOUR of NAND3_77 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_76 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_76;

architecture SYN_BEHAVIOUR of NAND3_76 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_75 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_75;

architecture SYN_BEHAVIOUR of NAND3_75 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_74 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_74;

architecture SYN_BEHAVIOUR of NAND3_74 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_73 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_73;

architecture SYN_BEHAVIOUR of NAND3_73 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_72 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_72;

architecture SYN_BEHAVIOUR of NAND3_72 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_71 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_71;

architecture SYN_BEHAVIOUR of NAND3_71 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_70 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_70;

architecture SYN_BEHAVIOUR of NAND3_70 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_69 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_69;

architecture SYN_BEHAVIOUR of NAND3_69 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_68 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_68;

architecture SYN_BEHAVIOUR of NAND3_68 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_67 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_67;

architecture SYN_BEHAVIOUR of NAND3_67 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_66 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_66;

architecture SYN_BEHAVIOUR of NAND3_66 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_65 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_65;

architecture SYN_BEHAVIOUR of NAND3_65 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_64 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_64;

architecture SYN_BEHAVIOUR of NAND3_64 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_63 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_63;

architecture SYN_BEHAVIOUR of NAND3_63 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_62 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_62;

architecture SYN_BEHAVIOUR of NAND3_62 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_61 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_61;

architecture SYN_BEHAVIOUR of NAND3_61 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_60 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_60;

architecture SYN_BEHAVIOUR of NAND3_60 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_59 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_59;

architecture SYN_BEHAVIOUR of NAND3_59 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_58 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_58;

architecture SYN_BEHAVIOUR of NAND3_58 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_57 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_57;

architecture SYN_BEHAVIOUR of NAND3_57 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_56 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_56;

architecture SYN_BEHAVIOUR of NAND3_56 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_55 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_55;

architecture SYN_BEHAVIOUR of NAND3_55 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_54 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_54;

architecture SYN_BEHAVIOUR of NAND3_54 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_53 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_53;

architecture SYN_BEHAVIOUR of NAND3_53 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_52 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_52;

architecture SYN_BEHAVIOUR of NAND3_52 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_51 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_51;

architecture SYN_BEHAVIOUR of NAND3_51 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_50 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_50;

architecture SYN_BEHAVIOUR of NAND3_50 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_49 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_49;

architecture SYN_BEHAVIOUR of NAND3_49 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_48 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_48;

architecture SYN_BEHAVIOUR of NAND3_48 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_47 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_47;

architecture SYN_BEHAVIOUR of NAND3_47 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_46 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_46;

architecture SYN_BEHAVIOUR of NAND3_46 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_45 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_45;

architecture SYN_BEHAVIOUR of NAND3_45 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_44 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_44;

architecture SYN_BEHAVIOUR of NAND3_44 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_43 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_43;

architecture SYN_BEHAVIOUR of NAND3_43 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_42 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_42;

architecture SYN_BEHAVIOUR of NAND3_42 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_41 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_41;

architecture SYN_BEHAVIOUR of NAND3_41 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_40 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_40;

architecture SYN_BEHAVIOUR of NAND3_40 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_39 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_39;

architecture SYN_BEHAVIOUR of NAND3_39 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_38 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_38;

architecture SYN_BEHAVIOUR of NAND3_38 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_37 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_37;

architecture SYN_BEHAVIOUR of NAND3_37 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_36 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_36;

architecture SYN_BEHAVIOUR of NAND3_36 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_35 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_35;

architecture SYN_BEHAVIOUR of NAND3_35 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_34 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_34;

architecture SYN_BEHAVIOUR of NAND3_34 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_33 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_33;

architecture SYN_BEHAVIOUR of NAND3_33 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_32 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_32;

architecture SYN_BEHAVIOUR of NAND3_32 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_31 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_31;

architecture SYN_BEHAVIOUR of NAND3_31 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_30 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_30;

architecture SYN_BEHAVIOUR of NAND3_30 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_29 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_29;

architecture SYN_BEHAVIOUR of NAND3_29 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_28 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_28;

architecture SYN_BEHAVIOUR of NAND3_28 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_27 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_27;

architecture SYN_BEHAVIOUR of NAND3_27 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_26 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_26;

architecture SYN_BEHAVIOUR of NAND3_26 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_25 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_25;

architecture SYN_BEHAVIOUR of NAND3_25 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_24 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_24;

architecture SYN_BEHAVIOUR of NAND3_24 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_23 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_23;

architecture SYN_BEHAVIOUR of NAND3_23 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_22 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_22;

architecture SYN_BEHAVIOUR of NAND3_22 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_21 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_21;

architecture SYN_BEHAVIOUR of NAND3_21 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_20 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_20;

architecture SYN_BEHAVIOUR of NAND3_20 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_19 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_19;

architecture SYN_BEHAVIOUR of NAND3_19 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_18 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_18;

architecture SYN_BEHAVIOUR of NAND3_18 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_17 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_17;

architecture SYN_BEHAVIOUR of NAND3_17 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_16 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_16;

architecture SYN_BEHAVIOUR of NAND3_16 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_15 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_15;

architecture SYN_BEHAVIOUR of NAND3_15 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_14 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_14;

architecture SYN_BEHAVIOUR of NAND3_14 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_13 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_13;

architecture SYN_BEHAVIOUR of NAND3_13 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_12 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_12;

architecture SYN_BEHAVIOUR of NAND3_12 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_11 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_11;

architecture SYN_BEHAVIOUR of NAND3_11 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_10 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_10;

architecture SYN_BEHAVIOUR of NAND3_10 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_9 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_9;

architecture SYN_BEHAVIOUR of NAND3_9 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_8 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_8;

architecture SYN_BEHAVIOUR of NAND3_8 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_7 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_7;

architecture SYN_BEHAVIOUR of NAND3_7 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_6 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_6;

architecture SYN_BEHAVIOUR of NAND3_6 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_5 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_5;

architecture SYN_BEHAVIOUR of NAND3_5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_4 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_4;

architecture SYN_BEHAVIOUR of NAND3_4 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_3 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_3;

architecture SYN_BEHAVIOUR of NAND3_3 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_2 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_2;

architecture SYN_BEHAVIOUR of NAND3_2 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_1 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_1;

architecture SYN_BEHAVIOUR of NAND3_1 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT5_1 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_GENERIC_NBIT5_1;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT5_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U5 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_4;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_3;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n33, n34, n35 : std_logic;

begin
   
   U1 : BUF_X4 port map( A => n35, Z => Y(0));
   U2 : BUF_X4 port map( A => n34, Z => Y(1));
   U3 : BUF_X4 port map( A => n33, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U5 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U6 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U7 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U8 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U9 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U10 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U11 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U12 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U13 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U14 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U15 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U16 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U17 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U20 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U23 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U24 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U25 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U26 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U27 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U28 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U29 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U30 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U31 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U32 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U33 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => n33);
   U34 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => n34);
   U35 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_2;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_1;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT5_2 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 downto 
         0);  DATA_OUT : out std_logic_vector (4 downto 0));

end REG_GENERIC_NBIT5_2;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT5_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n14, CK => CLK, Q => DATA_OUT(4)
                           , QN => n13);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n15, CK => CLK, Q => DATA_OUT(3)
                           , QN => n12);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n16, CK => CLK, Q => DATA_OUT(2)
                           , QN => n11);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n17, CK => CLK, Q => DATA_OUT(1)
                           , QN => n10);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n18, CK => CLK, Q => DATA_OUT(0)
                           , QN => n9);
   U3 : OAI21_X1 port map( B1 => n13, B2 => n1, A => n2, ZN => n14);
   U4 : NAND2_X1 port map( A1 => DATA_IN(4), A2 => n3, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n12, B2 => n1, A => n4, ZN => n15);
   U6 : NAND2_X1 port map( A1 => DATA_IN(3), A2 => n3, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n11, B2 => n1, A => n5, ZN => n16);
   U8 : NAND2_X1 port map( A1 => DATA_IN(2), A2 => n3, ZN => n5);
   U9 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n6, ZN => n17);
   U10 : NAND2_X1 port map( A1 => DATA_IN(1), A2 => n3, ZN => n6);
   U11 : OAI21_X1 port map( B1 => n9, B2 => n1, A => n7, ZN => n18);
   U12 : NAND2_X1 port map( A1 => DATA_IN(0), A2 => n3, ZN => n7);
   U13 : AND2_X1 port map( A1 => RST, A2 => n1, ZN => n3);
   U14 : NAND2_X1 port map( A1 => n8, A2 => RST, ZN => n1);
   U15 : INV_X1 port map( A => EN, ZN => n8);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT5_1 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 downto 
         0);  DATA_OUT : out std_logic_vector (4 downto 0));

end REG_GENERIC_NBIT5_1;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n14, CK => CLK, Q => DATA_OUT(4)
                           , QN => n13);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n15, CK => CLK, Q => DATA_OUT(3)
                           , QN => n12);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n16, CK => CLK, Q => DATA_OUT(2)
                           , QN => n11);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n17, CK => CLK, Q => DATA_OUT(1)
                           , QN => n10);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n18, CK => CLK, Q => DATA_OUT(0)
                           , QN => n9);
   U3 : OAI21_X1 port map( B1 => n13, B2 => n1, A => n2, ZN => n14);
   U4 : NAND2_X1 port map( A1 => DATA_IN(4), A2 => n3, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n12, B2 => n1, A => n4, ZN => n15);
   U6 : NAND2_X1 port map( A1 => DATA_IN(3), A2 => n3, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n11, B2 => n1, A => n5, ZN => n16);
   U8 : NAND2_X1 port map( A1 => DATA_IN(2), A2 => n3, ZN => n5);
   U9 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n6, ZN => n17);
   U10 : NAND2_X1 port map( A1 => DATA_IN(1), A2 => n3, ZN => n6);
   U11 : OAI21_X1 port map( B1 => n9, B2 => n1, A => n7, ZN => n18);
   U12 : NAND2_X1 port map( A1 => DATA_IN(0), A2 => n3, ZN => n7);
   U13 : AND2_X1 port map( A1 => RST, A2 => n1, ZN => n3);
   U14 : NAND2_X1 port map( A1 => n8, A2 => RST, ZN => n1);
   U15 : INV_X1 port map( A => EN, ZN => n8);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_8 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_8;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_7 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_7;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_6 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_6;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_5 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_5;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_4 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_4;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_3 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_3;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n91, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n93, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n92, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n90, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n81, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n80, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n86, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n68, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(0), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(31), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(26), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(27), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(24), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(25), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(30), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(28), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(29), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(23), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(10), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(11), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(8), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(9), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(14), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(15), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(12), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(13), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(7), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(18), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(19), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(16), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(17), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(22), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(20), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(21), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(2), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(3), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(1), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(6), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(4), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(5), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_2 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_2;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_1 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_1;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BARREL_SHIFTER_N32 is

   port( CONF : in std_logic;  DATA1, DATA2 : in std_logic_vector (31 downto 0)
         ;  OUTPUT : out std_logic_vector (31 downto 0));

end BARREL_SHIFTER_N32;

architecture SYN_BEHAVIOR of BARREL_SHIFTER_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal COARSE_39_port, COARSE_38_port, COARSE_37_port, COARSE_36_port, 
      COARSE_35_port, COARSE_34_port, COARSE_33_port, COARSE_32_port, 
      COARSE_31_port, COARSE_30_port, COARSE_29_port, COARSE_28_port, 
      COARSE_27_port, COARSE_26_port, COARSE_25_port, COARSE_24_port, 
      COARSE_23_port, COARSE_22_port, COARSE_21_port, COARSE_20_port, 
      COARSE_19_port, COARSE_18_port, COARSE_17_port, COARSE_16_port, 
      COARSE_15_port, COARSE_14_port, COARSE_13_port, COARSE_12_port, 
      COARSE_11_port, COARSE_10_port, COARSE_9_port, COARSE_8_port, 
      COARSE_7_port, COARSE_6_port, COARSE_5_port, COARSE_4_port, COARSE_3_port
      , COARSE_2_port, COARSE_1_port, COARSE_0_port, SL_OUT_31_port, 
      SL_OUT_30_port, SL_OUT_29_port, SL_OUT_28_port, SL_OUT_27_port, 
      SL_OUT_26_port, SL_OUT_25_port, SL_OUT_24_port, SL_OUT_23_port, 
      SL_OUT_22_port, SL_OUT_21_port, SL_OUT_20_port, SL_OUT_19_port, 
      SL_OUT_18_port, SL_OUT_17_port, SL_OUT_16_port, SL_OUT_15_port, 
      SL_OUT_14_port, SL_OUT_13_port, SL_OUT_12_port, SL_OUT_11_port, 
      SL_OUT_10_port, SL_OUT_9_port, SL_OUT_8_port, SL_OUT_7_port, 
      SL_OUT_6_port, SL_OUT_5_port, SL_OUT_4_port, SL_OUT_3_port, SL_OUT_2_port
      , SL_OUT_1_port, SL_OUT_0_port, SR_OUT_31_port, SR_OUT_30_port, 
      SR_OUT_29_port, SR_OUT_28_port, SR_OUT_27_port, SR_OUT_26_port, 
      SR_OUT_25_port, SR_OUT_24_port, SR_OUT_23_port, SR_OUT_22_port, 
      SR_OUT_21_port, SR_OUT_20_port, SR_OUT_19_port, SR_OUT_18_port, 
      SR_OUT_17_port, SR_OUT_16_port, SR_OUT_15_port, SR_OUT_14_port, 
      SR_OUT_13_port, SR_OUT_12_port, SR_OUT_11_port, SR_OUT_10_port, 
      SR_OUT_9_port, SR_OUT_8_port, SR_OUT_7_port, SR_OUT_6_port, SR_OUT_5_port
      , SR_OUT_4_port, SR_OUT_3_port, SR_OUT_2_port, SR_OUT_1_port, 
      SR_OUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325 : std_logic;

begin
   
   U2 : NOR3_X2 port map( A1 => n294, A2 => n241, A3 => n295, ZN => n255);
   U3 : NOR3_X4 port map( A1 => n241, A2 => DATA2(3), A3 => n294, ZN => n248);
   U4 : NOR3_X2 port map( A1 => n294, A2 => CONF, A3 => n295, ZN => n273);
   U5 : NAND3_X2 port map( A1 => n295, A2 => n294, A3 => CONF, ZN => n242);
   U6 : INV_X2 port map( A => CONF, ZN => n241);
   U7 : NOR3_X4 port map( A1 => CONF, A2 => DATA2(3), A3 => n294, ZN => n274);
   U8 : NOR3_X4 port map( A1 => CONF, A2 => DATA2(4), A3 => n295, ZN => n296);
   U9 : NOR3_X4 port map( A1 => DATA2(3), A2 => DATA2(4), A3 => CONF, ZN => 
                           n247);
   U10 : INV_X1 port map( A => COARSE_5_port, ZN => n162);
   U11 : INV_X1 port map( A => COARSE_4_port, ZN => n156);
   U12 : INV_X1 port map( A => COARSE_34_port, ZN => n146);
   U13 : INV_X1 port map( A => COARSE_35_port, ZN => n152);
   U14 : INV_X1 port map( A => n133, ZN => n164);
   U15 : INV_X1 port map( A => n12, ZN => n175);
   U16 : INV_X1 port map( A => n73, ZN => n209);
   U17 : INV_X1 port map( A => n69, ZN => n158);
   U18 : INV_X1 port map( A => COARSE_25_port, ZN => n145);
   U19 : INV_X1 port map( A => COARSE_24_port, ZN => n140);
   U20 : INV_X1 port map( A => COARSE_26_port, ZN => n150);
   U21 : INV_X1 port map( A => COARSE_27_port, ZN => n155);
   U22 : INV_X1 port map( A => COARSE_28_port, ZN => n161);
   U23 : INV_X1 port map( A => COARSE_29_port, ZN => n167);
   U24 : INV_X1 port map( A => COARSE_30_port, ZN => n196);
   U25 : INV_X1 port map( A => COARSE_31_port, ZN => n232);
   U26 : INV_X1 port map( A => COARSE_6_port, ZN => n168);
   U27 : INV_X1 port map( A => COARSE_7_port, ZN => n205);
   U28 : INV_X1 port map( A => COARSE_8_port, ZN => n137);
   U29 : INV_X1 port map( A => COARSE_9_port, ZN => n141);
   U30 : INV_X1 port map( A => COARSE_10_port, ZN => n149);
   U31 : INV_X1 port map( A => COARSE_11_port, ZN => n154);
   U32 : INV_X1 port map( A => COARSE_12_port, ZN => n160);
   U33 : INV_X1 port map( A => COARSE_13_port, ZN => n166);
   U34 : INV_X1 port map( A => COARSE_14_port, ZN => n187);
   U35 : INV_X1 port map( A => COARSE_15_port, ZN => n223);
   U36 : INV_X1 port map( A => COARSE_16_port, ZN => n139);
   U37 : INV_X1 port map( A => COARSE_17_port, ZN => n144);
   U38 : INV_X1 port map( A => COARSE_18_port, ZN => n148);
   U39 : INV_X1 port map( A => COARSE_19_port, ZN => n153);
   U40 : INV_X1 port map( A => COARSE_20_port, ZN => n159);
   U41 : INV_X1 port map( A => COARSE_21_port, ZN => n165);
   U42 : INV_X1 port map( A => COARSE_22_port, ZN => n178);
   U43 : INV_X1 port map( A => COARSE_23_port, ZN => n214);
   U44 : INV_X1 port map( A => COARSE_2_port, ZN => n147);
   U45 : INV_X1 port map( A => COARSE_3_port, ZN => n151);
   U46 : INV_X1 port map( A => COARSE_33_port, ZN => n142);
   U47 : INV_X1 port map( A => COARSE_32_port, ZN => n138);
   U48 : INV_X1 port map( A => COARSE_37_port, ZN => n163);
   U49 : INV_X1 port map( A => COARSE_36_port, ZN => n157);
   U50 : INV_X1 port map( A => n11, ZN => n212);
   U51 : INV_X1 port map( A => COARSE_1_port, ZN => n143);
   U52 : INV_X1 port map( A => n76, ZN => n171);
   U53 : INV_X1 port map( A => n14, ZN => n174);
   U54 : INV_X1 port map( A => n78, ZN => n208);
   U55 : INV_X1 port map( A => n16, ZN => n213);
   U56 : INV_X1 port map( A => n80, ZN => n169);
   U57 : INV_X1 port map( A => n18, ZN => n172);
   U58 : INV_X1 port map( A => n82, ZN => n206);
   U59 : INV_X1 port map( A => n20, ZN => n210);
   U60 : INV_X1 port map( A => n84, ZN => n170);
   U61 : INV_X1 port map( A => n22, ZN => n173);
   U62 : INV_X1 port map( A => n86, ZN => n207);
   U63 : INV_X1 port map( A => n24, ZN => n211);
   U64 : INV_X1 port map( A => n88, ZN => n190);
   U65 : INV_X1 port map( A => n26, ZN => n194);
   U66 : INV_X1 port map( A => n90, ZN => n226);
   U67 : INV_X1 port map( A => n28, ZN => n230);
   U68 : INV_X1 port map( A => n92, ZN => n191);
   U69 : INV_X1 port map( A => n30, ZN => n195);
   U70 : INV_X1 port map( A => n94, ZN => n227);
   U71 : INV_X1 port map( A => n32, ZN => n231);
   U72 : INV_X1 port map( A => n96, ZN => n188);
   U73 : INV_X1 port map( A => n34, ZN => n192);
   U74 : INV_X1 port map( A => n98, ZN => n224);
   U75 : INV_X1 port map( A => n36, ZN => n228);
   U76 : INV_X1 port map( A => n100, ZN => n189);
   U77 : INV_X1 port map( A => n38, ZN => n193);
   U78 : INV_X1 port map( A => n102, ZN => n225);
   U79 : INV_X1 port map( A => n40, ZN => n229);
   U80 : INV_X1 port map( A => n104, ZN => n181);
   U81 : INV_X1 port map( A => n42, ZN => n185);
   U82 : INV_X1 port map( A => n106, ZN => n217);
   U83 : INV_X1 port map( A => n44, ZN => n221);
   U84 : INV_X1 port map( A => n108, ZN => n182);
   U85 : INV_X1 port map( A => n46, ZN => n186);
   U86 : INV_X1 port map( A => n110, ZN => n218);
   U87 : INV_X1 port map( A => n48, ZN => n222);
   U88 : INV_X1 port map( A => n112, ZN => n179);
   U89 : INV_X1 port map( A => n50, ZN => n183);
   U90 : INV_X1 port map( A => n114, ZN => n215);
   U91 : INV_X1 port map( A => n52, ZN => n219);
   U92 : INV_X1 port map( A => n116, ZN => n180);
   U93 : INV_X1 port map( A => n54, ZN => n184);
   U94 : INV_X1 port map( A => n118, ZN => n216);
   U95 : INV_X1 port map( A => n56, ZN => n220);
   U96 : INV_X1 port map( A => n120, ZN => n199);
   U97 : INV_X1 port map( A => n58, ZN => n203);
   U98 : INV_X1 port map( A => n122, ZN => n235);
   U99 : INV_X1 port map( A => n60, ZN => n239);
   U100 : INV_X1 port map( A => n124, ZN => n200);
   U101 : INV_X1 port map( A => n62, ZN => n204);
   U102 : INV_X1 port map( A => n126, ZN => n236);
   U103 : INV_X1 port map( A => n64, ZN => n240);
   U104 : INV_X1 port map( A => n128, ZN => n197);
   U105 : INV_X1 port map( A => n66, ZN => n201);
   U106 : INV_X1 port map( A => n130, ZN => n233);
   U107 : INV_X1 port map( A => n68, ZN => n237);
   U108 : INV_X1 port map( A => n132, ZN => n198);
   U109 : INV_X1 port map( A => n70, ZN => n202);
   U110 : INV_X1 port map( A => n134, ZN => n234);
   U111 : INV_X1 port map( A => n72, ZN => n238);
   U112 : INV_X1 port map( A => n136, ZN => n177);
   U113 : INV_X1 port map( A => COARSE_38_port, ZN => n176);
   U114 : MUX2_X1 port map( A => COARSE_0_port, B => COARSE_4_port, S => 
                           DATA2(2), Z => n1);
   U115 : MUX2_X1 port map( A => n1, B => n175, S => DATA2(1), Z => n2);
   U116 : MUX2_X1 port map( A => n2, B => n212, S => DATA2(0), Z => 
                           SR_OUT_0_port);
   U117 : MUX2_X1 port map( A => n212, B => n174, S => DATA2(0), Z => 
                           SR_OUT_1_port);
   U118 : MUX2_X1 port map( A => n174, B => n213, S => DATA2(0), Z => 
                           SR_OUT_2_port);
   U119 : MUX2_X1 port map( A => n213, B => n172, S => DATA2(0), Z => 
                           SR_OUT_3_port);
   U120 : MUX2_X1 port map( A => n172, B => n210, S => DATA2(0), Z => 
                           SR_OUT_4_port);
   U121 : MUX2_X1 port map( A => n210, B => n173, S => DATA2(0), Z => 
                           SR_OUT_5_port);
   U122 : MUX2_X1 port map( A => n173, B => n211, S => DATA2(0), Z => 
                           SR_OUT_6_port);
   U123 : MUX2_X1 port map( A => n211, B => n194, S => DATA2(0), Z => 
                           SR_OUT_7_port);
   U124 : MUX2_X1 port map( A => n194, B => n230, S => DATA2(0), Z => 
                           SR_OUT_8_port);
   U125 : MUX2_X1 port map( A => n230, B => n195, S => DATA2(0), Z => 
                           SR_OUT_9_port);
   U126 : MUX2_X1 port map( A => n195, B => n231, S => DATA2(0), Z => 
                           SR_OUT_10_port);
   U127 : MUX2_X1 port map( A => n231, B => n192, S => DATA2(0), Z => 
                           SR_OUT_11_port);
   U128 : MUX2_X1 port map( A => n192, B => n228, S => DATA2(0), Z => 
                           SR_OUT_12_port);
   U129 : MUX2_X1 port map( A => n228, B => n193, S => DATA2(0), Z => 
                           SR_OUT_13_port);
   U130 : MUX2_X1 port map( A => n193, B => n229, S => DATA2(0), Z => 
                           SR_OUT_14_port);
   U131 : MUX2_X1 port map( A => n229, B => n185, S => DATA2(0), Z => 
                           SR_OUT_15_port);
   U132 : MUX2_X1 port map( A => n185, B => n221, S => DATA2(0), Z => 
                           SR_OUT_16_port);
   U133 : MUX2_X1 port map( A => n221, B => n186, S => DATA2(0), Z => 
                           SR_OUT_17_port);
   U134 : MUX2_X1 port map( A => n186, B => n222, S => DATA2(0), Z => 
                           SR_OUT_18_port);
   U135 : MUX2_X1 port map( A => n222, B => n183, S => DATA2(0), Z => 
                           SR_OUT_19_port);
   U136 : MUX2_X1 port map( A => n183, B => n219, S => DATA2(0), Z => 
                           SR_OUT_20_port);
   U137 : MUX2_X1 port map( A => n219, B => n184, S => DATA2(0), Z => 
                           SR_OUT_21_port);
   U138 : MUX2_X1 port map( A => n184, B => n220, S => DATA2(0), Z => 
                           SR_OUT_22_port);
   U139 : MUX2_X1 port map( A => n220, B => n203, S => DATA2(0), Z => 
                           SR_OUT_23_port);
   U140 : MUX2_X1 port map( A => n203, B => n239, S => DATA2(0), Z => 
                           SR_OUT_24_port);
   U141 : MUX2_X1 port map( A => n239, B => n204, S => DATA2(0), Z => 
                           SR_OUT_25_port);
   U142 : MUX2_X1 port map( A => n204, B => n240, S => DATA2(0), Z => 
                           SR_OUT_26_port);
   U143 : MUX2_X1 port map( A => n240, B => n201, S => DATA2(0), Z => 
                           SR_OUT_27_port);
   U144 : MUX2_X1 port map( A => n201, B => n237, S => DATA2(0), Z => 
                           SR_OUT_28_port);
   U145 : MUX2_X1 port map( A => n237, B => n202, S => DATA2(0), Z => 
                           SR_OUT_29_port);
   U146 : MUX2_X1 port map( A => n202, B => n238, S => DATA2(0), Z => 
                           SR_OUT_30_port);
   U147 : MUX2_X1 port map( A => COARSE_34_port, B => COARSE_38_port, S => 
                           DATA2(2), Z => n3);
   U148 : MUX2_X1 port map( A => n158, B => n3, S => DATA2(1), Z => n4);
   U149 : MUX2_X1 port map( A => n238, B => n4, S => DATA2(0), Z => 
                           SR_OUT_31_port);
   U150 : MUX2_X1 port map( A => COARSE_5_port, B => COARSE_1_port, S => 
                           DATA2(2), Z => n5);
   U151 : MUX2_X1 port map( A => n209, B => n5, S => DATA2(1), Z => n6);
   U152 : MUX2_X1 port map( A => n171, B => n6, S => DATA2(0), Z => 
                           SL_OUT_0_port);
   U153 : MUX2_X1 port map( A => n208, B => n171, S => DATA2(0), Z => 
                           SL_OUT_1_port);
   U154 : MUX2_X1 port map( A => n169, B => n208, S => DATA2(0), Z => 
                           SL_OUT_2_port);
   U155 : MUX2_X1 port map( A => n206, B => n169, S => DATA2(0), Z => 
                           SL_OUT_3_port);
   U156 : MUX2_X1 port map( A => n170, B => n206, S => DATA2(0), Z => 
                           SL_OUT_4_port);
   U157 : MUX2_X1 port map( A => n207, B => n170, S => DATA2(0), Z => 
                           SL_OUT_5_port);
   U158 : MUX2_X1 port map( A => n190, B => n207, S => DATA2(0), Z => 
                           SL_OUT_6_port);
   U159 : MUX2_X1 port map( A => n226, B => n190, S => DATA2(0), Z => 
                           SL_OUT_7_port);
   U160 : MUX2_X1 port map( A => n191, B => n226, S => DATA2(0), Z => 
                           SL_OUT_8_port);
   U161 : MUX2_X1 port map( A => n227, B => n191, S => DATA2(0), Z => 
                           SL_OUT_9_port);
   U162 : MUX2_X1 port map( A => n188, B => n227, S => DATA2(0), Z => 
                           SL_OUT_10_port);
   U163 : MUX2_X1 port map( A => n224, B => n188, S => DATA2(0), Z => 
                           SL_OUT_11_port);
   U164 : MUX2_X1 port map( A => n189, B => n224, S => DATA2(0), Z => 
                           SL_OUT_12_port);
   U165 : MUX2_X1 port map( A => n225, B => n189, S => DATA2(0), Z => 
                           SL_OUT_13_port);
   U166 : MUX2_X1 port map( A => n181, B => n225, S => DATA2(0), Z => 
                           SL_OUT_14_port);
   U167 : MUX2_X1 port map( A => n217, B => n181, S => DATA2(0), Z => 
                           SL_OUT_15_port);
   U168 : MUX2_X1 port map( A => n182, B => n217, S => DATA2(0), Z => 
                           SL_OUT_16_port);
   U169 : MUX2_X1 port map( A => n218, B => n182, S => DATA2(0), Z => 
                           SL_OUT_17_port);
   U170 : MUX2_X1 port map( A => n179, B => n218, S => DATA2(0), Z => 
                           SL_OUT_18_port);
   U171 : MUX2_X1 port map( A => n215, B => n179, S => DATA2(0), Z => 
                           SL_OUT_19_port);
   U172 : MUX2_X1 port map( A => n180, B => n215, S => DATA2(0), Z => 
                           SL_OUT_20_port);
   U173 : MUX2_X1 port map( A => n216, B => n180, S => DATA2(0), Z => 
                           SL_OUT_21_port);
   U174 : MUX2_X1 port map( A => n199, B => n216, S => DATA2(0), Z => 
                           SL_OUT_22_port);
   U175 : MUX2_X1 port map( A => n235, B => n199, S => DATA2(0), Z => 
                           SL_OUT_23_port);
   U176 : MUX2_X1 port map( A => n200, B => n235, S => DATA2(0), Z => 
                           SL_OUT_24_port);
   U177 : MUX2_X1 port map( A => n236, B => n200, S => DATA2(0), Z => 
                           SL_OUT_25_port);
   U178 : MUX2_X1 port map( A => n197, B => n236, S => DATA2(0), Z => 
                           SL_OUT_26_port);
   U179 : MUX2_X1 port map( A => n233, B => n197, S => DATA2(0), Z => 
                           SL_OUT_27_port);
   U180 : MUX2_X1 port map( A => n198, B => n233, S => DATA2(0), Z => 
                           SL_OUT_28_port);
   U181 : MUX2_X1 port map( A => n234, B => n198, S => DATA2(0), Z => 
                           SL_OUT_29_port);
   U182 : MUX2_X1 port map( A => n177, B => n234, S => DATA2(0), Z => 
                           SL_OUT_30_port);
   U183 : MUX2_X1 port map( A => COARSE_39_port, B => COARSE_35_port, S => 
                           DATA2(2), Z => n7);
   U184 : MUX2_X1 port map( A => n7, B => n164, S => DATA2(1), Z => n8);
   U185 : MUX2_X1 port map( A => n8, B => n177, S => DATA2(0), Z => 
                           SL_OUT_31_port);
   U186 : MUX2_X1 port map( A => n151, B => n205, S => DATA2(2), Z => n9);
   U187 : MUX2_X1 port map( A => n143, B => n162, S => DATA2(2), Z => n10);
   U188 : MUX2_X1 port map( A => n10, B => n9, S => DATA2(1), Z => n11);
   U189 : MUX2_X1 port map( A => n147, B => n168, S => DATA2(2), Z => n12);
   U190 : MUX2_X1 port map( A => n156, B => n137, S => DATA2(2), Z => n13);
   U191 : MUX2_X1 port map( A => n12, B => n13, S => DATA2(1), Z => n14);
   U192 : MUX2_X1 port map( A => n162, B => n141, S => DATA2(2), Z => n15);
   U193 : MUX2_X1 port map( A => n9, B => n15, S => DATA2(1), Z => n16);
   U194 : MUX2_X1 port map( A => n168, B => n149, S => DATA2(2), Z => n17);
   U195 : MUX2_X1 port map( A => n13, B => n17, S => DATA2(1), Z => n18);
   U196 : MUX2_X1 port map( A => n205, B => n154, S => DATA2(2), Z => n19);
   U197 : MUX2_X1 port map( A => n15, B => n19, S => DATA2(1), Z => n20);
   U198 : MUX2_X1 port map( A => n137, B => n160, S => DATA2(2), Z => n21);
   U199 : MUX2_X1 port map( A => n17, B => n21, S => DATA2(1), Z => n22);
   U200 : MUX2_X1 port map( A => n141, B => n166, S => DATA2(2), Z => n23);
   U201 : MUX2_X1 port map( A => n19, B => n23, S => DATA2(1), Z => n24);
   U202 : MUX2_X1 port map( A => n149, B => n187, S => DATA2(2), Z => n25);
   U203 : MUX2_X1 port map( A => n21, B => n25, S => DATA2(1), Z => n26);
   U204 : MUX2_X1 port map( A => n154, B => n223, S => DATA2(2), Z => n27);
   U205 : MUX2_X1 port map( A => n23, B => n27, S => DATA2(1), Z => n28);
   U206 : MUX2_X1 port map( A => n160, B => n139, S => DATA2(2), Z => n29);
   U207 : MUX2_X1 port map( A => n25, B => n29, S => DATA2(1), Z => n30);
   U208 : MUX2_X1 port map( A => n166, B => n144, S => DATA2(2), Z => n31);
   U209 : MUX2_X1 port map( A => n27, B => n31, S => DATA2(1), Z => n32);
   U210 : MUX2_X1 port map( A => n187, B => n148, S => DATA2(2), Z => n33);
   U211 : MUX2_X1 port map( A => n29, B => n33, S => DATA2(1), Z => n34);
   U212 : MUX2_X1 port map( A => n223, B => n153, S => DATA2(2), Z => n35);
   U213 : MUX2_X1 port map( A => n31, B => n35, S => DATA2(1), Z => n36);
   U214 : MUX2_X1 port map( A => n139, B => n159, S => DATA2(2), Z => n37);
   U215 : MUX2_X1 port map( A => n33, B => n37, S => DATA2(1), Z => n38);
   U216 : MUX2_X1 port map( A => n144, B => n165, S => DATA2(2), Z => n39);
   U217 : MUX2_X1 port map( A => n35, B => n39, S => DATA2(1), Z => n40);
   U218 : MUX2_X1 port map( A => n148, B => n178, S => DATA2(2), Z => n41);
   U219 : MUX2_X1 port map( A => n37, B => n41, S => DATA2(1), Z => n42);
   U220 : MUX2_X1 port map( A => n153, B => n214, S => DATA2(2), Z => n43);
   U221 : MUX2_X1 port map( A => n39, B => n43, S => DATA2(1), Z => n44);
   U222 : MUX2_X1 port map( A => n159, B => n140, S => DATA2(2), Z => n45);
   U223 : MUX2_X1 port map( A => n41, B => n45, S => DATA2(1), Z => n46);
   U224 : MUX2_X1 port map( A => n165, B => n145, S => DATA2(2), Z => n47);
   U225 : MUX2_X1 port map( A => n43, B => n47, S => DATA2(1), Z => n48);
   U226 : MUX2_X1 port map( A => n178, B => n150, S => DATA2(2), Z => n49);
   U227 : MUX2_X1 port map( A => n45, B => n49, S => DATA2(1), Z => n50);
   U228 : MUX2_X1 port map( A => n214, B => n155, S => DATA2(2), Z => n51);
   U229 : MUX2_X1 port map( A => n47, B => n51, S => DATA2(1), Z => n52);
   U230 : MUX2_X1 port map( A => n140, B => n161, S => DATA2(2), Z => n53);
   U231 : MUX2_X1 port map( A => n49, B => n53, S => DATA2(1), Z => n54);
   U232 : MUX2_X1 port map( A => n145, B => n167, S => DATA2(2), Z => n55);
   U233 : MUX2_X1 port map( A => n51, B => n55, S => DATA2(1), Z => n56);
   U234 : MUX2_X1 port map( A => n150, B => n196, S => DATA2(2), Z => n57);
   U235 : MUX2_X1 port map( A => n53, B => n57, S => DATA2(1), Z => n58);
   U236 : MUX2_X1 port map( A => n155, B => n232, S => DATA2(2), Z => n59);
   U237 : MUX2_X1 port map( A => n55, B => n59, S => DATA2(1), Z => n60);
   U238 : MUX2_X1 port map( A => n161, B => n138, S => DATA2(2), Z => n61);
   U239 : MUX2_X1 port map( A => n57, B => n61, S => DATA2(1), Z => n62);
   U240 : MUX2_X1 port map( A => n167, B => n142, S => DATA2(2), Z => n63);
   U241 : MUX2_X1 port map( A => n59, B => n63, S => DATA2(1), Z => n64);
   U242 : MUX2_X1 port map( A => n196, B => n146, S => DATA2(2), Z => n65);
   U243 : MUX2_X1 port map( A => n61, B => n65, S => DATA2(1), Z => n66);
   U244 : MUX2_X1 port map( A => n232, B => n152, S => DATA2(2), Z => n67);
   U245 : MUX2_X1 port map( A => n63, B => n67, S => DATA2(1), Z => n68);
   U246 : MUX2_X1 port map( A => n138, B => n157, S => DATA2(2), Z => n69);
   U247 : MUX2_X1 port map( A => n65, B => n69, S => DATA2(1), Z => n70);
   U248 : MUX2_X1 port map( A => n142, B => n163, S => DATA2(2), Z => n71);
   U249 : MUX2_X1 port map( A => n67, B => n71, S => DATA2(1), Z => n72);
   U250 : MUX2_X1 port map( A => n205, B => n151, S => DATA2(2), Z => n73);
   U251 : MUX2_X1 port map( A => n168, B => n147, S => DATA2(2), Z => n74);
   U252 : MUX2_X1 port map( A => n137, B => n156, S => DATA2(2), Z => n75);
   U253 : MUX2_X1 port map( A => n75, B => n74, S => DATA2(1), Z => n76);
   U254 : MUX2_X1 port map( A => n141, B => n162, S => DATA2(2), Z => n77);
   U255 : MUX2_X1 port map( A => n77, B => n73, S => DATA2(1), Z => n78);
   U256 : MUX2_X1 port map( A => n149, B => n168, S => DATA2(2), Z => n79);
   U257 : MUX2_X1 port map( A => n79, B => n75, S => DATA2(1), Z => n80);
   U258 : MUX2_X1 port map( A => n154, B => n205, S => DATA2(2), Z => n81);
   U259 : MUX2_X1 port map( A => n81, B => n77, S => DATA2(1), Z => n82);
   U260 : MUX2_X1 port map( A => n160, B => n137, S => DATA2(2), Z => n83);
   U261 : MUX2_X1 port map( A => n83, B => n79, S => DATA2(1), Z => n84);
   U262 : MUX2_X1 port map( A => n166, B => n141, S => DATA2(2), Z => n85);
   U263 : MUX2_X1 port map( A => n85, B => n81, S => DATA2(1), Z => n86);
   U264 : MUX2_X1 port map( A => n187, B => n149, S => DATA2(2), Z => n87);
   U265 : MUX2_X1 port map( A => n87, B => n83, S => DATA2(1), Z => n88);
   U266 : MUX2_X1 port map( A => n223, B => n154, S => DATA2(2), Z => n89);
   U267 : MUX2_X1 port map( A => n89, B => n85, S => DATA2(1), Z => n90);
   U268 : MUX2_X1 port map( A => n139, B => n160, S => DATA2(2), Z => n91);
   U269 : MUX2_X1 port map( A => n91, B => n87, S => DATA2(1), Z => n92);
   U270 : MUX2_X1 port map( A => n144, B => n166, S => DATA2(2), Z => n93);
   U271 : MUX2_X1 port map( A => n93, B => n89, S => DATA2(1), Z => n94);
   U272 : MUX2_X1 port map( A => n148, B => n187, S => DATA2(2), Z => n95);
   U273 : MUX2_X1 port map( A => n95, B => n91, S => DATA2(1), Z => n96);
   U274 : MUX2_X1 port map( A => n153, B => n223, S => DATA2(2), Z => n97);
   U275 : MUX2_X1 port map( A => n97, B => n93, S => DATA2(1), Z => n98);
   U276 : MUX2_X1 port map( A => n159, B => n139, S => DATA2(2), Z => n99);
   U277 : MUX2_X1 port map( A => n99, B => n95, S => DATA2(1), Z => n100);
   U278 : MUX2_X1 port map( A => n165, B => n144, S => DATA2(2), Z => n101);
   U279 : MUX2_X1 port map( A => n101, B => n97, S => DATA2(1), Z => n102);
   U280 : MUX2_X1 port map( A => n178, B => n148, S => DATA2(2), Z => n103);
   U281 : MUX2_X1 port map( A => n103, B => n99, S => DATA2(1), Z => n104);
   U282 : MUX2_X1 port map( A => n214, B => n153, S => DATA2(2), Z => n105);
   U283 : MUX2_X1 port map( A => n105, B => n101, S => DATA2(1), Z => n106);
   U284 : MUX2_X1 port map( A => n140, B => n159, S => DATA2(2), Z => n107);
   U285 : MUX2_X1 port map( A => n107, B => n103, S => DATA2(1), Z => n108);
   U286 : MUX2_X1 port map( A => n145, B => n165, S => DATA2(2), Z => n109);
   U287 : MUX2_X1 port map( A => n109, B => n105, S => DATA2(1), Z => n110);
   U288 : MUX2_X1 port map( A => n150, B => n178, S => DATA2(2), Z => n111);
   U289 : MUX2_X1 port map( A => n111, B => n107, S => DATA2(1), Z => n112);
   U290 : MUX2_X1 port map( A => n155, B => n214, S => DATA2(2), Z => n113);
   U291 : MUX2_X1 port map( A => n113, B => n109, S => DATA2(1), Z => n114);
   U292 : MUX2_X1 port map( A => n161, B => n140, S => DATA2(2), Z => n115);
   U293 : MUX2_X1 port map( A => n115, B => n111, S => DATA2(1), Z => n116);
   U294 : MUX2_X1 port map( A => n167, B => n145, S => DATA2(2), Z => n117);
   U295 : MUX2_X1 port map( A => n117, B => n113, S => DATA2(1), Z => n118);
   U296 : MUX2_X1 port map( A => n196, B => n150, S => DATA2(2), Z => n119);
   U297 : MUX2_X1 port map( A => n119, B => n115, S => DATA2(1), Z => n120);
   U298 : MUX2_X1 port map( A => n232, B => n155, S => DATA2(2), Z => n121);
   U299 : MUX2_X1 port map( A => n121, B => n117, S => DATA2(1), Z => n122);
   U300 : MUX2_X1 port map( A => n138, B => n161, S => DATA2(2), Z => n123);
   U301 : MUX2_X1 port map( A => n123, B => n119, S => DATA2(1), Z => n124);
   U302 : MUX2_X1 port map( A => n142, B => n167, S => DATA2(2), Z => n125);
   U303 : MUX2_X1 port map( A => n125, B => n121, S => DATA2(1), Z => n126);
   U304 : MUX2_X1 port map( A => n146, B => n196, S => DATA2(2), Z => n127);
   U305 : MUX2_X1 port map( A => n127, B => n123, S => DATA2(1), Z => n128);
   U306 : MUX2_X1 port map( A => n152, B => n232, S => DATA2(2), Z => n129);
   U307 : MUX2_X1 port map( A => n129, B => n125, S => DATA2(1), Z => n130);
   U308 : MUX2_X1 port map( A => n157, B => n138, S => DATA2(2), Z => n131);
   U309 : MUX2_X1 port map( A => n131, B => n127, S => DATA2(1), Z => n132);
   U310 : MUX2_X1 port map( A => n163, B => n142, S => DATA2(2), Z => n133);
   U311 : MUX2_X1 port map( A => n133, B => n129, S => DATA2(1), Z => n134);
   U312 : MUX2_X1 port map( A => n176, B => n146, S => DATA2(2), Z => n135);
   U313 : MUX2_X1 port map( A => n135, B => n131, S => DATA2(1), Z => n136);
   U314 : MUX2_X1 port map( A => SR_OUT_26_port, B => SL_OUT_26_port, S => n241
                           , Z => OUTPUT(26));
   U315 : MUX2_X1 port map( A => SR_OUT_27_port, B => SL_OUT_27_port, S => n241
                           , Z => OUTPUT(27));
   U316 : MUX2_X1 port map( A => SR_OUT_24_port, B => SL_OUT_24_port, S => n241
                           , Z => OUTPUT(24));
   U317 : MUX2_X1 port map( A => SR_OUT_25_port, B => SL_OUT_25_port, S => n241
                           , Z => OUTPUT(25));
   U318 : MUX2_X1 port map( A => SR_OUT_30_port, B => SL_OUT_30_port, S => n241
                           , Z => OUTPUT(30));
   U319 : MUX2_X1 port map( A => SR_OUT_31_port, B => SL_OUT_31_port, S => n241
                           , Z => OUTPUT(31));
   U320 : MUX2_X1 port map( A => SR_OUT_28_port, B => SL_OUT_28_port, S => n241
                           , Z => OUTPUT(28));
   U321 : MUX2_X1 port map( A => SR_OUT_29_port, B => SL_OUT_29_port, S => n241
                           , Z => OUTPUT(29));
   U322 : MUX2_X1 port map( A => SR_OUT_23_port, B => SL_OUT_23_port, S => n241
                           , Z => OUTPUT(23));
   U323 : MUX2_X1 port map( A => SR_OUT_10_port, B => SL_OUT_10_port, S => n241
                           , Z => OUTPUT(10));
   U324 : MUX2_X1 port map( A => SR_OUT_11_port, B => SL_OUT_11_port, S => n241
                           , Z => OUTPUT(11));
   U325 : MUX2_X1 port map( A => SR_OUT_8_port, B => SL_OUT_8_port, S => n241, 
                           Z => OUTPUT(8));
   U326 : MUX2_X1 port map( A => SR_OUT_9_port, B => SL_OUT_9_port, S => n241, 
                           Z => OUTPUT(9));
   U327 : MUX2_X1 port map( A => SR_OUT_14_port, B => SL_OUT_14_port, S => n241
                           , Z => OUTPUT(14));
   U328 : MUX2_X1 port map( A => SR_OUT_15_port, B => SL_OUT_15_port, S => n241
                           , Z => OUTPUT(15));
   U329 : MUX2_X1 port map( A => SR_OUT_12_port, B => SL_OUT_12_port, S => n241
                           , Z => OUTPUT(12));
   U330 : MUX2_X1 port map( A => SR_OUT_13_port, B => SL_OUT_13_port, S => n241
                           , Z => OUTPUT(13));
   U331 : MUX2_X1 port map( A => SR_OUT_7_port, B => SL_OUT_7_port, S => n241, 
                           Z => OUTPUT(7));
   U332 : MUX2_X1 port map( A => SR_OUT_18_port, B => SL_OUT_18_port, S => n241
                           , Z => OUTPUT(18));
   U333 : MUX2_X1 port map( A => SR_OUT_19_port, B => SL_OUT_19_port, S => n241
                           , Z => OUTPUT(19));
   U334 : MUX2_X1 port map( A => SR_OUT_16_port, B => SL_OUT_16_port, S => n241
                           , Z => OUTPUT(16));
   U335 : MUX2_X1 port map( A => SR_OUT_17_port, B => SL_OUT_17_port, S => n241
                           , Z => OUTPUT(17));
   U336 : MUX2_X1 port map( A => SR_OUT_22_port, B => SL_OUT_22_port, S => n241
                           , Z => OUTPUT(22));
   U337 : MUX2_X1 port map( A => SR_OUT_20_port, B => SL_OUT_20_port, S => n241
                           , Z => OUTPUT(20));
   U338 : MUX2_X1 port map( A => SR_OUT_21_port, B => SL_OUT_21_port, S => n241
                           , Z => OUTPUT(21));
   U339 : MUX2_X1 port map( A => SR_OUT_2_port, B => SL_OUT_2_port, S => n241, 
                           Z => OUTPUT(2));
   U340 : MUX2_X1 port map( A => SR_OUT_3_port, B => SL_OUT_3_port, S => n241, 
                           Z => OUTPUT(3));
   U341 : MUX2_X1 port map( A => SR_OUT_0_port, B => SL_OUT_0_port, S => n241, 
                           Z => OUTPUT(0));
   U342 : MUX2_X1 port map( A => SR_OUT_1_port, B => SL_OUT_1_port, S => n241, 
                           Z => OUTPUT(1));
   U343 : MUX2_X1 port map( A => SR_OUT_6_port, B => SL_OUT_6_port, S => n241, 
                           Z => OUTPUT(6));
   U344 : MUX2_X1 port map( A => SR_OUT_4_port, B => SL_OUT_4_port, S => n241, 
                           Z => OUTPUT(4));
   U345 : MUX2_X1 port map( A => SR_OUT_5_port, B => SL_OUT_5_port, S => n241, 
                           Z => OUTPUT(5));
   U346 : OAI221_X1 port map( B1 => n242, B2 => n243, C1 => n244, C2 => n245, A
                           => n246, ZN => COARSE_9_port);
   U347 : AOI22_X1 port map( A1 => DATA1(1), A2 => n247, B1 => DATA1(25), B2 =>
                           n248, ZN => n246);
   U348 : OAI221_X1 port map( B1 => n242, B2 => n249, C1 => n244, C2 => n250, A
                           => n251, ZN => COARSE_8_port);
   U349 : AOI22_X1 port map( A1 => DATA1(0), A2 => n247, B1 => DATA1(24), B2 =>
                           n248, ZN => n251);
   U350 : OAI221_X1 port map( B1 => n242, B2 => n252, C1 => n244, C2 => n253, A
                           => n254, ZN => COARSE_7_port);
   U351 : AOI22_X1 port map( A1 => DATA1(23), A2 => n248, B1 => DATA1(31), B2 
                           => n255, ZN => n254);
   U352 : INV_X1 port map( A => DATA1(7), ZN => n252);
   U353 : OAI221_X1 port map( B1 => n242, B2 => n256, C1 => n244, C2 => n257, A
                           => n258, ZN => COARSE_6_port);
   U354 : AOI22_X1 port map( A1 => DATA1(22), A2 => n248, B1 => DATA1(30), B2 
                           => n255, ZN => n258);
   U355 : INV_X1 port map( A => DATA1(6), ZN => n256);
   U356 : OAI221_X1 port map( B1 => n242, B2 => n259, C1 => n244, C2 => n260, A
                           => n261, ZN => COARSE_5_port);
   U357 : AOI22_X1 port map( A1 => DATA1(21), A2 => n248, B1 => DATA1(29), B2 
                           => n255, ZN => n261);
   U358 : INV_X1 port map( A => DATA1(5), ZN => n259);
   U359 : OAI221_X1 port map( B1 => n242, B2 => n262, C1 => n244, C2 => n263, A
                           => n264, ZN => COARSE_4_port);
   U360 : AOI22_X1 port map( A1 => DATA1(20), A2 => n248, B1 => DATA1(28), B2 
                           => n255, ZN => n264);
   U361 : INV_X1 port map( A => DATA1(4), ZN => n262);
   U362 : OAI221_X1 port map( B1 => n242, B2 => n265, C1 => n244, C2 => n266, A
                           => n267, ZN => COARSE_3_port);
   U363 : AOI22_X1 port map( A1 => DATA1(19), A2 => n248, B1 => DATA1(27), B2 
                           => n255, ZN => n267);
   U364 : INV_X1 port map( A => DATA1(3), ZN => n265);
   U365 : OAI221_X1 port map( B1 => n268, B2 => n269, C1 => n270, C2 => n271, A
                           => n272, ZN => COARSE_39_port);
   U366 : AOI22_X1 port map( A1 => n273, A2 => DATA1(7), B1 => n274, B2 => 
                           DATA1(15), ZN => n272);
   U367 : OAI221_X1 port map( B1 => n275, B2 => n269, C1 => n270, C2 => n276, A
                           => n277, ZN => COARSE_38_port);
   U368 : AOI22_X1 port map( A1 => n273, A2 => DATA1(6), B1 => n274, B2 => 
                           DATA1(14), ZN => n277);
   U369 : OAI221_X1 port map( B1 => n278, B2 => n269, C1 => n270, C2 => n279, A
                           => n280, ZN => COARSE_37_port);
   U370 : AOI22_X1 port map( A1 => n273, A2 => DATA1(5), B1 => n274, B2 => 
                           DATA1(13), ZN => n280);
   U371 : OAI221_X1 port map( B1 => n281, B2 => n269, C1 => n270, C2 => n282, A
                           => n283, ZN => COARSE_36_port);
   U372 : AOI22_X1 port map( A1 => n273, A2 => DATA1(4), B1 => n274, B2 => 
                           DATA1(12), ZN => n283);
   U373 : OAI221_X1 port map( B1 => n284, B2 => n269, C1 => n270, C2 => n285, A
                           => n286, ZN => COARSE_35_port);
   U374 : AOI22_X1 port map( A1 => n273, A2 => DATA1(3), B1 => n274, B2 => 
                           DATA1(11), ZN => n286);
   U375 : OAI221_X1 port map( B1 => n269, B2 => n287, C1 => n270, C2 => n288, A
                           => n289, ZN => COARSE_34_port);
   U376 : AOI22_X1 port map( A1 => DATA1(2), A2 => n273, B1 => DATA1(10), B2 =>
                           n274, ZN => n289);
   U377 : OAI221_X1 port map( B1 => n245, B2 => n269, C1 => n270, C2 => n290, A
                           => n291, ZN => COARSE_33_port);
   U378 : AOI22_X1 port map( A1 => n273, A2 => DATA1(1), B1 => n274, B2 => 
                           DATA1(9), ZN => n291);
   U379 : OAI221_X1 port map( B1 => n250, B2 => n269, C1 => n270, C2 => n292, A
                           => n293, ZN => COARSE_32_port);
   U380 : AOI22_X1 port map( A1 => n273, A2 => DATA1(0), B1 => n274, B2 => 
                           DATA1(8), ZN => n293);
   U381 : INV_X1 port map( A => n296, ZN => n269);
   U382 : OAI221_X1 port map( B1 => n270, B2 => n268, C1 => n242, C2 => n271, A
                           => n297, ZN => COARSE_31_port);
   U383 : AOI22_X1 port map( A1 => n274, A2 => DATA1(7), B1 => n296, B2 => 
                           DATA1(15), ZN => n297);
   U384 : OAI221_X1 port map( B1 => n270, B2 => n275, C1 => n242, C2 => n276, A
                           => n298, ZN => COARSE_30_port);
   U385 : AOI22_X1 port map( A1 => n274, A2 => DATA1(6), B1 => n296, B2 => 
                           DATA1(14), ZN => n298);
   U386 : OAI221_X1 port map( B1 => n242, B2 => n299, C1 => n244, C2 => n300, A
                           => n301, ZN => COARSE_2_port);
   U387 : AOI22_X1 port map( A1 => DATA1(18), A2 => n248, B1 => DATA1(26), B2 
                           => n255, ZN => n301);
   U388 : INV_X1 port map( A => DATA1(2), ZN => n299);
   U389 : OAI221_X1 port map( B1 => n270, B2 => n278, C1 => n242, C2 => n279, A
                           => n302, ZN => COARSE_29_port);
   U390 : AOI22_X1 port map( A1 => n274, A2 => DATA1(5), B1 => n296, B2 => 
                           DATA1(13), ZN => n302);
   U391 : OAI221_X1 port map( B1 => n270, B2 => n281, C1 => n242, C2 => n282, A
                           => n303, ZN => COARSE_28_port);
   U392 : AOI22_X1 port map( A1 => n274, A2 => DATA1(4), B1 => n296, B2 => 
                           DATA1(12), ZN => n303);
   U393 : OAI221_X1 port map( B1 => n270, B2 => n284, C1 => n242, C2 => n285, A
                           => n304, ZN => COARSE_27_port);
   U394 : AOI22_X1 port map( A1 => n274, A2 => DATA1(3), B1 => n296, B2 => 
                           DATA1(11), ZN => n304);
   U395 : OAI221_X1 port map( B1 => n270, B2 => n287, C1 => n242, C2 => n288, A
                           => n305, ZN => COARSE_26_port);
   U396 : AOI22_X1 port map( A1 => DATA1(2), A2 => n274, B1 => DATA1(10), B2 =>
                           n296, ZN => n305);
   U397 : OAI221_X1 port map( B1 => n270, B2 => n245, C1 => n290, C2 => n242, A
                           => n306, ZN => COARSE_25_port);
   U398 : AOI22_X1 port map( A1 => n274, A2 => DATA1(1), B1 => n296, B2 => 
                           DATA1(9), ZN => n306);
   U399 : OAI221_X1 port map( B1 => n270, B2 => n250, C1 => n242, C2 => n292, A
                           => n307, ZN => COARSE_24_port);
   U400 : AOI22_X1 port map( A1 => n274, A2 => DATA1(0), B1 => n296, B2 => 
                           DATA1(8), ZN => n307);
   U401 : INV_X1 port map( A => n247, ZN => n270);
   U402 : OAI221_X1 port map( B1 => n242, B2 => n268, C1 => n244, C2 => n271, A
                           => n308, ZN => COARSE_23_port);
   U403 : AOI22_X1 port map( A1 => n296, A2 => DATA1(7), B1 => DATA1(15), B2 =>
                           n247, ZN => n308);
   U404 : INV_X1 port map( A => DATA1(31), ZN => n271);
   U405 : OAI221_X1 port map( B1 => n242, B2 => n275, C1 => n244, C2 => n276, A
                           => n309, ZN => COARSE_22_port);
   U406 : AOI22_X1 port map( A1 => n296, A2 => DATA1(6), B1 => DATA1(14), B2 =>
                           n247, ZN => n309);
   U407 : INV_X1 port map( A => DATA1(30), ZN => n276);
   U408 : OAI221_X1 port map( B1 => n242, B2 => n278, C1 => n244, C2 => n279, A
                           => n310, ZN => COARSE_21_port);
   U409 : AOI22_X1 port map( A1 => n296, A2 => DATA1(5), B1 => DATA1(13), B2 =>
                           n247, ZN => n310);
   U410 : INV_X1 port map( A => DATA1(29), ZN => n279);
   U411 : OAI221_X1 port map( B1 => n242, B2 => n281, C1 => n244, C2 => n282, A
                           => n311, ZN => COARSE_20_port);
   U412 : AOI22_X1 port map( A1 => n296, A2 => DATA1(4), B1 => DATA1(12), B2 =>
                           n247, ZN => n311);
   U413 : INV_X1 port map( A => DATA1(28), ZN => n282);
   U414 : OAI221_X1 port map( B1 => n312, B2 => n242, C1 => n243, C2 => n244, A
                           => n313, ZN => COARSE_1_port);
   U415 : AOI22_X1 port map( A1 => DATA1(17), A2 => n248, B1 => n255, B2 => 
                           DATA1(25), ZN => n313);
   U416 : INV_X1 port map( A => DATA1(9), ZN => n243);
   U417 : INV_X1 port map( A => DATA1(1), ZN => n312);
   U418 : OAI221_X1 port map( B1 => n242, B2 => n284, C1 => n244, C2 => n285, A
                           => n314, ZN => COARSE_19_port);
   U419 : AOI22_X1 port map( A1 => n296, A2 => DATA1(3), B1 => DATA1(11), B2 =>
                           n247, ZN => n314);
   U420 : INV_X1 port map( A => DATA1(27), ZN => n285);
   U421 : OAI221_X1 port map( B1 => n242, B2 => n287, C1 => n244, C2 => n288, A
                           => n315, ZN => COARSE_18_port);
   U422 : AOI22_X1 port map( A1 => DATA1(2), A2 => n296, B1 => DATA1(10), B2 =>
                           n247, ZN => n315);
   U423 : INV_X1 port map( A => DATA1(26), ZN => n288);
   U424 : OAI221_X1 port map( B1 => n242, B2 => n245, C1 => n290, C2 => n244, A
                           => n316, ZN => COARSE_17_port);
   U425 : AOI22_X1 port map( A1 => n296, A2 => DATA1(1), B1 => DATA1(9), B2 => 
                           n247, ZN => n316);
   U426 : INV_X1 port map( A => DATA1(25), ZN => n290);
   U427 : INV_X1 port map( A => DATA1(17), ZN => n245);
   U428 : OAI221_X1 port map( B1 => n242, B2 => n250, C1 => n244, C2 => n292, A
                           => n317, ZN => COARSE_16_port);
   U429 : AOI22_X1 port map( A1 => n296, A2 => DATA1(0), B1 => DATA1(8), B2 => 
                           n247, ZN => n317);
   U430 : INV_X1 port map( A => DATA1(24), ZN => n292);
   U431 : INV_X1 port map( A => DATA1(16), ZN => n250);
   U432 : OAI221_X1 port map( B1 => n242, B2 => n253, C1 => n244, C2 => n268, A
                           => n318, ZN => COARSE_15_port);
   U433 : AOI22_X1 port map( A1 => DATA1(7), A2 => n247, B1 => DATA1(31), B2 =>
                           n248, ZN => n318);
   U434 : INV_X1 port map( A => DATA1(23), ZN => n268);
   U435 : INV_X1 port map( A => DATA1(15), ZN => n253);
   U436 : OAI221_X1 port map( B1 => n242, B2 => n257, C1 => n244, C2 => n275, A
                           => n319, ZN => COARSE_14_port);
   U437 : AOI22_X1 port map( A1 => DATA1(6), A2 => n247, B1 => DATA1(30), B2 =>
                           n248, ZN => n319);
   U438 : INV_X1 port map( A => DATA1(22), ZN => n275);
   U439 : INV_X1 port map( A => DATA1(14), ZN => n257);
   U440 : OAI221_X1 port map( B1 => n242, B2 => n260, C1 => n244, C2 => n278, A
                           => n320, ZN => COARSE_13_port);
   U441 : AOI22_X1 port map( A1 => DATA1(5), A2 => n247, B1 => DATA1(29), B2 =>
                           n248, ZN => n320);
   U442 : INV_X1 port map( A => DATA1(21), ZN => n278);
   U443 : INV_X1 port map( A => DATA1(13), ZN => n260);
   U444 : OAI221_X1 port map( B1 => n242, B2 => n263, C1 => n244, C2 => n281, A
                           => n321, ZN => COARSE_12_port);
   U445 : AOI22_X1 port map( A1 => DATA1(4), A2 => n247, B1 => DATA1(28), B2 =>
                           n248, ZN => n321);
   U446 : INV_X1 port map( A => DATA1(20), ZN => n281);
   U447 : INV_X1 port map( A => DATA1(12), ZN => n263);
   U448 : OAI221_X1 port map( B1 => n242, B2 => n266, C1 => n244, C2 => n284, A
                           => n322, ZN => COARSE_11_port);
   U449 : AOI22_X1 port map( A1 => DATA1(3), A2 => n247, B1 => DATA1(27), B2 =>
                           n248, ZN => n322);
   U450 : INV_X1 port map( A => DATA1(19), ZN => n284);
   U451 : INV_X1 port map( A => DATA1(11), ZN => n266);
   U452 : OAI221_X1 port map( B1 => n242, B2 => n300, C1 => n244, C2 => n287, A
                           => n323, ZN => COARSE_10_port);
   U453 : AOI22_X1 port map( A1 => DATA1(2), A2 => n247, B1 => DATA1(26), B2 =>
                           n248, ZN => n323);
   U454 : INV_X1 port map( A => DATA1(18), ZN => n287);
   U455 : INV_X1 port map( A => DATA1(10), ZN => n300);
   U456 : OAI221_X1 port map( B1 => n242, B2 => n324, C1 => n244, C2 => n249, A
                           => n325, ZN => COARSE_0_port);
   U457 : AOI22_X1 port map( A1 => DATA1(16), A2 => n248, B1 => n255, B2 => 
                           DATA1(24), ZN => n325);
   U458 : INV_X1 port map( A => DATA1(8), ZN => n249);
   U459 : NAND3_X1 port map( A1 => CONF, A2 => n294, A3 => DATA2(3), ZN => n244
                           );
   U460 : INV_X1 port map( A => DATA1(0), ZN => n324);
   U461 : INV_X1 port map( A => DATA2(4), ZN => n294);
   U462 : INV_X1 port map( A => DATA2(3), ZN => n295);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND4_0 is

   port( A, B, C, D : in std_logic;  Y : out std_logic);

end NAND4_0;

architecture SYN_BEHAVIOUR of NAND4_0 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => D, A2 => C, A3 => B, A4 => A, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity NAND3_0 is

   port( A, B, C : in std_logic;  Y : out std_logic);

end NAND3_0;

architecture SYN_BEHAVIOUR of NAND3_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => B, A2 => A, A3 => C, ZN => Y);

end SYN_BEHAVIOUR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32 is

   port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
         downto 0));

end ALU_N32;

architecture SYN_BEHAVIOR of ALU_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ALU_N32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component ALU_N32_DW01_addsub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (31 downto 0);  CO : out 
            std_logic);
   end component;
   
   component BARREL_SHIFTER_N32
      port( CONF : in std_logic;  DATA1, DATA2 : in std_logic_vector (31 downto
            0);  OUTPUT : out std_logic_vector (31 downto 0));
   end component;
   
   component NAND4_1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_2
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_3
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_4
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_5
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_6
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_7
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_8
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_9
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_10
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_11
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_12
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_13
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_14
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_15
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_16
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_17
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_18
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_19
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_20
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_21
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_22
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_23
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_24
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_25
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_26
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_27
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_28
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_29
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_30
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_31
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND4_0
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_2
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_3
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_4
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_5
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_6
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_7
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_8
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_9
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_10
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_11
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_12
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_13
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_14
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_15
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_16
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_17
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_18
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_19
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_20
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_21
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_22
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_23
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_24
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_25
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_26
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_27
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_28
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_29
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_30
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_31
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_32
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_33
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_34
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_35
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_36
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_37
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_38
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_39
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_40
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_41
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_42
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_43
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_44
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_45
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_46
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_47
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_48
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_49
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_50
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_51
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_52
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_53
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_54
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_55
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_56
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_57
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_58
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_59
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_60
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_61
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_62
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_63
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_64
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_65
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_66
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_67
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_68
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_69
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_70
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_71
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_72
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_73
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_74
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_75
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_76
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_77
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_78
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_79
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_80
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_81
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_82
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_83
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_84
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_85
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_86
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_87
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_88
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_89
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_90
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_91
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_92
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_93
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_94
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_95
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_96
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_97
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_98
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_99
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_100
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_101
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_102
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_103
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_104
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_105
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_106
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_107
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_108
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_109
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_110
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_111
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_112
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_113
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_114
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_115
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_116
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_117
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_118
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_119
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_120
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_121
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_122
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_123
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_124
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_125
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_126
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_127
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3_0
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89,
      N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
      N104, N105, N106, N107, N108, N109, N110, Y_LOGIC_31_port, 
      Y_LOGIC_30_port, Y_LOGIC_29_port, Y_LOGIC_28_port, Y_LOGIC_27_port, 
      Y_LOGIC_26_port, Y_LOGIC_25_port, Y_LOGIC_24_port, Y_LOGIC_23_port, 
      Y_LOGIC_22_port, Y_LOGIC_21_port, Y_LOGIC_20_port, Y_LOGIC_19_port, 
      Y_LOGIC_18_port, Y_LOGIC_17_port, Y_LOGIC_16_port, Y_LOGIC_15_port, 
      Y_LOGIC_14_port, Y_LOGIC_13_port, Y_LOGIC_12_port, Y_LOGIC_11_port, 
      Y_LOGIC_10_port, Y_LOGIC_9_port, Y_LOGIC_8_port, Y_LOGIC_7_port, 
      Y_LOGIC_6_port, Y_LOGIC_5_port, Y_LOGIC_4_port, Y_LOGIC_3_port, 
      Y_LOGIC_2_port, Y_LOGIC_1_port, Y_LOGIC_0_port, N111, N112, N113, 
      OUT_SHIFTER_31_port, OUT_SHIFTER_30_port, OUT_SHIFTER_29_port, 
      OUT_SHIFTER_28_port, OUT_SHIFTER_27_port, OUT_SHIFTER_26_port, 
      OUT_SHIFTER_25_port, OUT_SHIFTER_24_port, OUT_SHIFTER_23_port, 
      OUT_SHIFTER_22_port, OUT_SHIFTER_21_port, OUT_SHIFTER_20_port, 
      OUT_SHIFTER_19_port, OUT_SHIFTER_18_port, OUT_SHIFTER_17_port, 
      OUT_SHIFTER_16_port, OUT_SHIFTER_15_port, OUT_SHIFTER_14_port, 
      OUT_SHIFTER_13_port, OUT_SHIFTER_12_port, OUT_SHIFTER_11_port, 
      OUT_SHIFTER_10_port, OUT_SHIFTER_9_port, OUT_SHIFTER_8_port, 
      OUT_SHIFTER_7_port, OUT_SHIFTER_6_port, OUT_SHIFTER_5_port, 
      OUT_SHIFTER_4_port, OUT_SHIFTER_3_port, OUT_SHIFTER_2_port, 
      OUT_SHIFTER_1_port, OUT_SHIFTER_0_port, S_3_port, S_2_port, L0_31_port, 
      L0_30_port, L0_29_port, L0_28_port, L0_27_port, L0_26_port, L0_25_port, 
      L0_24_port, L0_23_port, L0_22_port, L0_21_port, L0_20_port, L0_19_port, 
      L0_18_port, L0_17_port, L0_16_port, L0_15_port, L0_14_port, L0_13_port, 
      L0_12_port, L0_11_port, L0_10_port, L0_9_port, L0_8_port, L0_7_port, 
      L0_6_port, L0_5_port, L0_4_port, L0_3_port, L0_2_port, L0_1_port, 
      L0_0_port, L1_31_port, L1_30_port, L1_29_port, L1_28_port, L1_27_port, 
      L1_26_port, L1_25_port, L1_24_port, L1_23_port, L1_22_port, L1_21_port, 
      L1_20_port, L1_19_port, L1_18_port, L1_17_port, L1_16_port, L1_15_port, 
      L1_14_port, L1_13_port, L1_12_port, L1_11_port, L1_10_port, L1_9_port, 
      L1_8_port, L1_7_port, L1_6_port, L1_5_port, L1_4_port, L1_3_port, 
      L1_2_port, L1_1_port, L1_0_port, L2_31_port, L2_30_port, L2_29_port, 
      L2_28_port, L2_27_port, L2_26_port, L2_25_port, L2_24_port, L2_23_port, 
      L2_22_port, L2_21_port, L2_20_port, L2_19_port, L2_18_port, L2_17_port, 
      L2_16_port, L2_15_port, L2_14_port, L2_13_port, L2_12_port, L2_11_port, 
      L2_10_port, L2_9_port, L2_8_port, L2_7_port, L2_6_port, L2_5_port, 
      L2_4_port, L2_3_port, L2_2_port, L2_1_port, L2_0_port, L3_31_port, 
      L3_30_port, L3_29_port, L3_28_port, L3_27_port, L3_26_port, L3_25_port, 
      L3_24_port, L3_23_port, L3_22_port, L3_21_port, L3_20_port, L3_19_port, 
      L3_18_port, L3_17_port, L3_16_port, L3_15_port, L3_14_port, L3_13_port, 
      L3_12_port, L3_11_port, L3_10_port, L3_9_port, L3_8_port, L3_7_port, 
      L3_6_port, L3_5_port, L3_4_port, L3_3_port, L3_2_port, L3_1_port, 
      L3_0_port, U2_U1_Z_0, U2_U2_Z_0, n12, n160, n1, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n84_port, n85_port, n86_port, n87_port, n88_port, n89_port, n90_port, 
      n91_port, n92_port, n93_port, n94_port, n95_port, n96_port, n97_port, 
      n98_port, n99_port, n100_port, n101_port, n102_port, n103_port, n104_port
      , n105_port, n106_port, n107_port, n108_port, n109_port, n110_port, 
      n111_port, n112_port, n113_port, n114, n115, n116, n117, n118, n119, n120
      , n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n_1040, n_1041, n_1042, n_1043 : std_logic;

begin
   
   X_Logic0_port <= '0';
   n12 <= '0';
   NAND31I_1 : NAND3_0 port map( A => n115, B => n147, C => X_Logic0_port, Y =>
                           L0_0_port);
   NAND31I_2 : NAND3_127 port map( A => n114, B => n146, C => X_Logic0_port, Y 
                           => L0_1_port);
   NAND31I_3 : NAND3_126 port map( A => n113_port, B => n145, C => 
                           X_Logic0_port, Y => L0_2_port);
   NAND31I_4 : NAND3_125 port map( A => n112_port, B => n144, C => 
                           X_Logic0_port, Y => L0_3_port);
   NAND31I_5 : NAND3_124 port map( A => n111_port, B => n143, C => 
                           X_Logic0_port, Y => L0_4_port);
   NAND31I_6 : NAND3_123 port map( A => n110_port, B => n142, C => 
                           X_Logic0_port, Y => L0_5_port);
   NAND31I_7 : NAND3_122 port map( A => n109_port, B => n141, C => 
                           X_Logic0_port, Y => L0_6_port);
   NAND31I_8 : NAND3_121 port map( A => n108_port, B => n140, C => 
                           X_Logic0_port, Y => L0_7_port);
   NAND31I_9 : NAND3_120 port map( A => n107_port, B => n139, C => 
                           X_Logic0_port, Y => L0_8_port);
   NAND31I_10 : NAND3_119 port map( A => n106_port, B => n138, C => 
                           X_Logic0_port, Y => L0_9_port);
   NAND31I_11 : NAND3_118 port map( A => n105_port, B => n137, C => 
                           X_Logic0_port, Y => L0_10_port);
   NAND31I_12 : NAND3_117 port map( A => n104_port, B => n136, C => 
                           X_Logic0_port, Y => L0_11_port);
   NAND31I_13 : NAND3_116 port map( A => n103_port, B => n135, C => 
                           X_Logic0_port, Y => L0_12_port);
   NAND31I_14 : NAND3_115 port map( A => n102_port, B => n134, C => 
                           X_Logic0_port, Y => L0_13_port);
   NAND31I_15 : NAND3_114 port map( A => n101_port, B => n133, C => 
                           X_Logic0_port, Y => L0_14_port);
   NAND31I_16 : NAND3_113 port map( A => n100_port, B => n132, C => 
                           X_Logic0_port, Y => L0_15_port);
   NAND31I_17 : NAND3_112 port map( A => n99_port, B => n131, C => 
                           X_Logic0_port, Y => L0_16_port);
   NAND31I_18 : NAND3_111 port map( A => n98_port, B => n130, C => 
                           X_Logic0_port, Y => L0_17_port);
   NAND31I_19 : NAND3_110 port map( A => n97_port, B => n129, C => 
                           X_Logic0_port, Y => L0_18_port);
   NAND31I_20 : NAND3_109 port map( A => n96_port, B => n128, C => 
                           X_Logic0_port, Y => L0_19_port);
   NAND31I_21 : NAND3_108 port map( A => n95_port, B => n127, C => 
                           X_Logic0_port, Y => L0_20_port);
   NAND31I_22 : NAND3_107 port map( A => n94_port, B => n126, C => 
                           X_Logic0_port, Y => L0_21_port);
   NAND31I_23 : NAND3_106 port map( A => n93_port, B => n125, C => 
                           X_Logic0_port, Y => L0_22_port);
   NAND31I_24 : NAND3_105 port map( A => n92_port, B => n124, C => 
                           X_Logic0_port, Y => L0_23_port);
   NAND31I_25 : NAND3_104 port map( A => n91_port, B => n123, C => 
                           X_Logic0_port, Y => L0_24_port);
   NAND31I_26 : NAND3_103 port map( A => n90_port, B => n122, C => 
                           X_Logic0_port, Y => L0_25_port);
   NAND31I_27 : NAND3_102 port map( A => n89_port, B => n121, C => 
                           X_Logic0_port, Y => L0_26_port);
   NAND31I_28 : NAND3_101 port map( A => n88_port, B => n120, C => 
                           X_Logic0_port, Y => L0_27_port);
   NAND31I_29 : NAND3_100 port map( A => n87_port, B => n119, C => 
                           X_Logic0_port, Y => L0_28_port);
   NAND31I_30 : NAND3_99 port map( A => n86_port, B => n118, C => X_Logic0_port
                           , Y => L0_29_port);
   NAND31I_31 : NAND3_98 port map( A => n85_port, B => n117, C => X_Logic0_port
                           , Y => L0_30_port);
   NAND31I_32 : NAND3_97 port map( A => n84_port, B => n116, C => X_Logic0_port
                           , Y => L0_31_port);
   NAND31I_1_0 : NAND3_96 port map( A => n115, B => DATA2(0), C => S_2_port, Y 
                           => L1_0_port);
   NAND31I_2_0 : NAND3_95 port map( A => n114, B => DATA2(1), C => S_2_port, Y 
                           => L1_1_port);
   NAND31I_3_0 : NAND3_94 port map( A => n113_port, B => DATA2(2), C => 
                           S_2_port, Y => L1_2_port);
   NAND31I_4_0 : NAND3_93 port map( A => n112_port, B => DATA2(3), C => 
                           S_2_port, Y => L1_3_port);
   NAND31I_5_0 : NAND3_92 port map( A => n111_port, B => DATA2(4), C => 
                           S_2_port, Y => L1_4_port);
   NAND31I_6_0 : NAND3_91 port map( A => n110_port, B => DATA2(5), C => 
                           S_2_port, Y => L1_5_port);
   NAND31I_7_0 : NAND3_90 port map( A => n109_port, B => DATA2(6), C => 
                           S_2_port, Y => L1_6_port);
   NAND31I_8_0 : NAND3_89 port map( A => n108_port, B => DATA2(7), C => 
                           S_2_port, Y => L1_7_port);
   NAND31I_9_0 : NAND3_88 port map( A => n107_port, B => DATA2(8), C => 
                           S_2_port, Y => L1_8_port);
   NAND31I_10_0 : NAND3_87 port map( A => n106_port, B => DATA2(9), C => 
                           S_2_port, Y => L1_9_port);
   NAND31I_11_0 : NAND3_86 port map( A => n105_port, B => DATA2(10), C => 
                           S_2_port, Y => L1_10_port);
   NAND31I_12_0 : NAND3_85 port map( A => n104_port, B => DATA2(11), C => 
                           S_2_port, Y => L1_11_port);
   NAND31I_13_0 : NAND3_84 port map( A => n103_port, B => DATA2(12), C => 
                           S_2_port, Y => L1_12_port);
   NAND31I_14_0 : NAND3_83 port map( A => n102_port, B => DATA2(13), C => 
                           S_2_port, Y => L1_13_port);
   NAND31I_15_0 : NAND3_82 port map( A => n101_port, B => DATA2(14), C => 
                           S_2_port, Y => L1_14_port);
   NAND31I_16_0 : NAND3_81 port map( A => n100_port, B => DATA2(15), C => 
                           S_2_port, Y => L1_15_port);
   NAND31I_17_0 : NAND3_80 port map( A => n99_port, B => DATA2(16), C => 
                           S_2_port, Y => L1_16_port);
   NAND31I_18_0 : NAND3_79 port map( A => n98_port, B => DATA2(17), C => 
                           S_2_port, Y => L1_17_port);
   NAND31I_19_0 : NAND3_78 port map( A => n97_port, B => DATA2(18), C => 
                           S_2_port, Y => L1_18_port);
   NAND31I_20_0 : NAND3_77 port map( A => n96_port, B => DATA2(19), C => 
                           S_2_port, Y => L1_19_port);
   NAND31I_21_0 : NAND3_76 port map( A => n95_port, B => DATA2(20), C => 
                           S_2_port, Y => L1_20_port);
   NAND31I_22_0 : NAND3_75 port map( A => n94_port, B => DATA2(21), C => 
                           S_2_port, Y => L1_21_port);
   NAND31I_23_0 : NAND3_74 port map( A => n93_port, B => DATA2(22), C => 
                           S_2_port, Y => L1_22_port);
   NAND31I_24_0 : NAND3_73 port map( A => n92_port, B => DATA2(23), C => 
                           S_2_port, Y => L1_23_port);
   NAND31I_25_0 : NAND3_72 port map( A => n91_port, B => DATA2(24), C => 
                           S_2_port, Y => L1_24_port);
   NAND31I_26_0 : NAND3_71 port map( A => n90_port, B => DATA2(25), C => 
                           S_2_port, Y => L1_25_port);
   NAND31I_27_0 : NAND3_70 port map( A => n89_port, B => DATA2(26), C => 
                           S_2_port, Y => L1_26_port);
   NAND31I_28_0 : NAND3_69 port map( A => n88_port, B => DATA2(27), C => 
                           S_2_port, Y => L1_27_port);
   NAND31I_29_0 : NAND3_68 port map( A => n87_port, B => DATA2(28), C => 
                           S_2_port, Y => L1_28_port);
   NAND31I_30_0 : NAND3_67 port map( A => n86_port, B => DATA2(29), C => 
                           S_2_port, Y => L1_29_port);
   NAND31I_31_0 : NAND3_66 port map( A => n85_port, B => DATA2(30), C => 
                           S_2_port, Y => L1_30_port);
   NAND31I_32_0 : NAND3_65 port map( A => n84_port, B => DATA2(31), C => 
                           S_2_port, Y => L1_31_port);
   NAND31I_1_1 : NAND3_64 port map( A => DATA1(0), B => n147, C => S_2_port, Y 
                           => L2_0_port);
   NAND31I_2_1 : NAND3_63 port map( A => DATA1(1), B => n146, C => S_2_port, Y 
                           => L2_1_port);
   NAND31I_3_1 : NAND3_62 port map( A => DATA1(2), B => n145, C => S_2_port, Y 
                           => L2_2_port);
   NAND31I_4_1 : NAND3_61 port map( A => DATA1(3), B => n144, C => S_2_port, Y 
                           => L2_3_port);
   NAND31I_5_1 : NAND3_60 port map( A => DATA1(4), B => n143, C => S_2_port, Y 
                           => L2_4_port);
   NAND31I_6_1 : NAND3_59 port map( A => DATA1(5), B => n142, C => S_2_port, Y 
                           => L2_5_port);
   NAND31I_7_1 : NAND3_58 port map( A => DATA1(6), B => n141, C => S_2_port, Y 
                           => L2_6_port);
   NAND31I_8_1 : NAND3_57 port map( A => DATA1(7), B => n140, C => S_2_port, Y 
                           => L2_7_port);
   NAND31I_9_1 : NAND3_56 port map( A => DATA1(8), B => n139, C => S_2_port, Y 
                           => L2_8_port);
   NAND31I_10_1 : NAND3_55 port map( A => DATA1(9), B => n138, C => S_2_port, Y
                           => L2_9_port);
   NAND31I_11_1 : NAND3_54 port map( A => DATA1(10), B => n137, C => S_2_port, 
                           Y => L2_10_port);
   NAND31I_12_1 : NAND3_53 port map( A => DATA1(11), B => n136, C => S_2_port, 
                           Y => L2_11_port);
   NAND31I_13_1 : NAND3_52 port map( A => DATA1(12), B => n135, C => S_2_port, 
                           Y => L2_12_port);
   NAND31I_14_1 : NAND3_51 port map( A => DATA1(13), B => n134, C => S_2_port, 
                           Y => L2_13_port);
   NAND31I_15_1 : NAND3_50 port map( A => DATA1(14), B => n133, C => S_2_port, 
                           Y => L2_14_port);
   NAND31I_16_1 : NAND3_49 port map( A => DATA1(15), B => n132, C => S_2_port, 
                           Y => L2_15_port);
   NAND31I_17_1 : NAND3_48 port map( A => DATA1(16), B => n131, C => S_2_port, 
                           Y => L2_16_port);
   NAND31I_18_1 : NAND3_47 port map( A => DATA1(17), B => n130, C => S_2_port, 
                           Y => L2_17_port);
   NAND31I_19_1 : NAND3_46 port map( A => DATA1(18), B => n129, C => S_2_port, 
                           Y => L2_18_port);
   NAND31I_20_1 : NAND3_45 port map( A => DATA1(19), B => n128, C => S_2_port, 
                           Y => L2_19_port);
   NAND31I_21_1 : NAND3_44 port map( A => DATA1(20), B => n127, C => S_2_port, 
                           Y => L2_20_port);
   NAND31I_22_1 : NAND3_43 port map( A => DATA1(21), B => n126, C => S_2_port, 
                           Y => L2_21_port);
   NAND31I_23_1 : NAND3_42 port map( A => DATA1(22), B => n125, C => S_2_port, 
                           Y => L2_22_port);
   NAND31I_24_1 : NAND3_41 port map( A => DATA1(23), B => n124, C => S_2_port, 
                           Y => L2_23_port);
   NAND31I_25_1 : NAND3_40 port map( A => DATA1(24), B => n123, C => S_2_port, 
                           Y => L2_24_port);
   NAND31I_26_1 : NAND3_39 port map( A => DATA1(25), B => n122, C => S_2_port, 
                           Y => L2_25_port);
   NAND31I_27_1 : NAND3_38 port map( A => DATA1(26), B => n121, C => S_2_port, 
                           Y => L2_26_port);
   NAND31I_28_1 : NAND3_37 port map( A => DATA1(27), B => n120, C => S_2_port, 
                           Y => L2_27_port);
   NAND31I_29_1 : NAND3_36 port map( A => DATA1(28), B => n119, C => S_2_port, 
                           Y => L2_28_port);
   NAND31I_30_1 : NAND3_35 port map( A => DATA1(29), B => n118, C => S_2_port, 
                           Y => L2_29_port);
   NAND31I_31_1 : NAND3_34 port map( A => DATA1(30), B => n117, C => S_2_port, 
                           Y => L2_30_port);
   NAND31I_32_1 : NAND3_33 port map( A => DATA1(31), B => n116, C => S_2_port, 
                           Y => L2_31_port);
   NAND31I_1_2 : NAND3_32 port map( A => DATA1(0), B => DATA2(0), C => S_3_port
                           , Y => L3_0_port);
   NAND31I_2_2 : NAND3_31 port map( A => DATA1(1), B => DATA2(1), C => S_3_port
                           , Y => L3_1_port);
   NAND31I_3_2 : NAND3_30 port map( A => DATA1(2), B => DATA2(2), C => S_3_port
                           , Y => L3_2_port);
   NAND31I_4_2 : NAND3_29 port map( A => DATA1(3), B => DATA2(3), C => S_3_port
                           , Y => L3_3_port);
   NAND31I_5_2 : NAND3_28 port map( A => DATA1(4), B => DATA2(4), C => S_3_port
                           , Y => L3_4_port);
   NAND31I_6_2 : NAND3_27 port map( A => DATA1(5), B => DATA2(5), C => S_3_port
                           , Y => L3_5_port);
   NAND31I_7_2 : NAND3_26 port map( A => DATA1(6), B => DATA2(6), C => S_3_port
                           , Y => L3_6_port);
   NAND31I_8_2 : NAND3_25 port map( A => DATA1(7), B => DATA2(7), C => S_3_port
                           , Y => L3_7_port);
   NAND31I_9_2 : NAND3_24 port map( A => DATA1(8), B => DATA2(8), C => S_3_port
                           , Y => L3_8_port);
   NAND31I_10_2 : NAND3_23 port map( A => DATA1(9), B => DATA2(9), C => 
                           S_3_port, Y => L3_9_port);
   NAND31I_11_2 : NAND3_22 port map( A => DATA1(10), B => DATA2(10), C => 
                           S_3_port, Y => L3_10_port);
   NAND31I_12_2 : NAND3_21 port map( A => DATA1(11), B => DATA2(11), C => 
                           S_3_port, Y => L3_11_port);
   NAND31I_13_2 : NAND3_20 port map( A => DATA1(12), B => DATA2(12), C => 
                           S_3_port, Y => L3_12_port);
   NAND31I_14_2 : NAND3_19 port map( A => DATA1(13), B => DATA2(13), C => 
                           S_3_port, Y => L3_13_port);
   NAND31I_15_2 : NAND3_18 port map( A => DATA1(14), B => DATA2(14), C => 
                           S_3_port, Y => L3_14_port);
   NAND31I_16_2 : NAND3_17 port map( A => DATA1(15), B => DATA2(15), C => 
                           S_3_port, Y => L3_15_port);
   NAND31I_17_2 : NAND3_16 port map( A => DATA1(16), B => DATA2(16), C => 
                           S_3_port, Y => L3_16_port);
   NAND31I_18_2 : NAND3_15 port map( A => DATA1(17), B => DATA2(17), C => 
                           S_3_port, Y => L3_17_port);
   NAND31I_19_2 : NAND3_14 port map( A => DATA1(18), B => DATA2(18), C => 
                           S_3_port, Y => L3_18_port);
   NAND31I_20_2 : NAND3_13 port map( A => DATA1(19), B => DATA2(19), C => 
                           S_3_port, Y => L3_19_port);
   NAND31I_21_2 : NAND3_12 port map( A => DATA1(20), B => DATA2(20), C => 
                           S_3_port, Y => L3_20_port);
   NAND31I_22_2 : NAND3_11 port map( A => DATA1(21), B => DATA2(21), C => 
                           S_3_port, Y => L3_21_port);
   NAND31I_23_2 : NAND3_10 port map( A => DATA1(22), B => DATA2(22), C => 
                           S_3_port, Y => L3_22_port);
   NAND31I_24_2 : NAND3_9 port map( A => DATA1(23), B => DATA2(23), C => 
                           S_3_port, Y => L3_23_port);
   NAND31I_25_2 : NAND3_8 port map( A => DATA1(24), B => DATA2(24), C => 
                           S_3_port, Y => L3_24_port);
   NAND31I_26_2 : NAND3_7 port map( A => DATA1(25), B => DATA2(25), C => 
                           S_3_port, Y => L3_25_port);
   NAND31I_27_2 : NAND3_6 port map( A => DATA1(26), B => DATA2(26), C => 
                           S_3_port, Y => L3_26_port);
   NAND31I_28_2 : NAND3_5 port map( A => DATA1(27), B => DATA2(27), C => 
                           S_3_port, Y => L3_27_port);
   NAND31I_29_2 : NAND3_4 port map( A => DATA1(28), B => DATA2(28), C => 
                           S_3_port, Y => L3_28_port);
   NAND31I_30_2 : NAND3_3 port map( A => DATA1(29), B => DATA2(29), C => 
                           S_3_port, Y => L3_29_port);
   NAND31I_31_2 : NAND3_2 port map( A => DATA1(30), B => DATA2(30), C => 
                           S_3_port, Y => L3_30_port);
   NAND31I_32_2 : NAND3_1 port map( A => DATA1(31), B => DATA2(31), C => 
                           S_3_port, Y => L3_31_port);
   NAND41I_1 : NAND4_0 port map( A => L0_0_port, B => L1_0_port, C => L2_0_port
                           , D => L3_0_port, Y => Y_LOGIC_0_port);
   NAND41I_2 : NAND4_31 port map( A => L0_1_port, B => L1_1_port, C => 
                           L2_1_port, D => L3_1_port, Y => Y_LOGIC_1_port);
   NAND41I_3 : NAND4_30 port map( A => L0_2_port, B => L1_2_port, C => 
                           L2_2_port, D => L3_2_port, Y => Y_LOGIC_2_port);
   NAND41I_4 : NAND4_29 port map( A => L0_3_port, B => L1_3_port, C => 
                           L2_3_port, D => L3_3_port, Y => Y_LOGIC_3_port);
   NAND41I_5 : NAND4_28 port map( A => L0_4_port, B => L1_4_port, C => 
                           L2_4_port, D => L3_4_port, Y => Y_LOGIC_4_port);
   NAND41I_6 : NAND4_27 port map( A => L0_5_port, B => L1_5_port, C => 
                           L2_5_port, D => L3_5_port, Y => Y_LOGIC_5_port);
   NAND41I_7 : NAND4_26 port map( A => L0_6_port, B => L1_6_port, C => 
                           L2_6_port, D => L3_6_port, Y => Y_LOGIC_6_port);
   NAND41I_8 : NAND4_25 port map( A => L0_7_port, B => L1_7_port, C => 
                           L2_7_port, D => L3_7_port, Y => Y_LOGIC_7_port);
   NAND41I_9 : NAND4_24 port map( A => L0_8_port, B => L1_8_port, C => 
                           L2_8_port, D => L3_8_port, Y => Y_LOGIC_8_port);
   NAND41I_10 : NAND4_23 port map( A => L0_9_port, B => L1_9_port, C => 
                           L2_9_port, D => L3_9_port, Y => Y_LOGIC_9_port);
   NAND41I_11 : NAND4_22 port map( A => L0_10_port, B => L1_10_port, C => 
                           L2_10_port, D => L3_10_port, Y => Y_LOGIC_10_port);
   NAND41I_12 : NAND4_21 port map( A => L0_11_port, B => L1_11_port, C => 
                           L2_11_port, D => L3_11_port, Y => Y_LOGIC_11_port);
   NAND41I_13 : NAND4_20 port map( A => L0_12_port, B => L1_12_port, C => 
                           L2_12_port, D => L3_12_port, Y => Y_LOGIC_12_port);
   NAND41I_14 : NAND4_19 port map( A => L0_13_port, B => L1_13_port, C => 
                           L2_13_port, D => L3_13_port, Y => Y_LOGIC_13_port);
   NAND41I_15 : NAND4_18 port map( A => L0_14_port, B => L1_14_port, C => 
                           L2_14_port, D => L3_14_port, Y => Y_LOGIC_14_port);
   NAND41I_16 : NAND4_17 port map( A => L0_15_port, B => L1_15_port, C => 
                           L2_15_port, D => L3_15_port, Y => Y_LOGIC_15_port);
   NAND41I_17 : NAND4_16 port map( A => L0_16_port, B => L1_16_port, C => 
                           L2_16_port, D => L3_16_port, Y => Y_LOGIC_16_port);
   NAND41I_18 : NAND4_15 port map( A => L0_17_port, B => L1_17_port, C => 
                           L2_17_port, D => L3_17_port, Y => Y_LOGIC_17_port);
   NAND41I_19 : NAND4_14 port map( A => L0_18_port, B => L1_18_port, C => 
                           L2_18_port, D => L3_18_port, Y => Y_LOGIC_18_port);
   NAND41I_20 : NAND4_13 port map( A => L0_19_port, B => L1_19_port, C => 
                           L2_19_port, D => L3_19_port, Y => Y_LOGIC_19_port);
   NAND41I_21 : NAND4_12 port map( A => L0_20_port, B => L1_20_port, C => 
                           L2_20_port, D => L3_20_port, Y => Y_LOGIC_20_port);
   NAND41I_22 : NAND4_11 port map( A => L0_21_port, B => L1_21_port, C => 
                           L2_21_port, D => L3_21_port, Y => Y_LOGIC_21_port);
   NAND41I_23 : NAND4_10 port map( A => L0_22_port, B => L1_22_port, C => 
                           L2_22_port, D => L3_22_port, Y => Y_LOGIC_22_port);
   NAND41I_24 : NAND4_9 port map( A => L0_23_port, B => L1_23_port, C => 
                           L2_23_port, D => L3_23_port, Y => Y_LOGIC_23_port);
   NAND41I_25 : NAND4_8 port map( A => L0_24_port, B => L1_24_port, C => 
                           L2_24_port, D => L3_24_port, Y => Y_LOGIC_24_port);
   NAND41I_26 : NAND4_7 port map( A => L0_25_port, B => L1_25_port, C => 
                           L2_25_port, D => L3_25_port, Y => Y_LOGIC_25_port);
   NAND41I_27 : NAND4_6 port map( A => L0_26_port, B => L1_26_port, C => 
                           L2_26_port, D => L3_26_port, Y => Y_LOGIC_26_port);
   NAND41I_28 : NAND4_5 port map( A => L0_27_port, B => L1_27_port, C => 
                           L2_27_port, D => L3_27_port, Y => Y_LOGIC_27_port);
   NAND41I_29 : NAND4_4 port map( A => L0_28_port, B => L1_28_port, C => 
                           L2_28_port, D => L3_28_port, Y => Y_LOGIC_28_port);
   NAND41I_30 : NAND4_3 port map( A => L0_29_port, B => L1_29_port, C => 
                           L2_29_port, D => L3_29_port, Y => Y_LOGIC_29_port);
   NAND41I_31 : NAND4_2 port map( A => L0_30_port, B => L1_30_port, C => 
                           L2_30_port, D => L3_30_port, Y => Y_LOGIC_30_port);
   NAND41I_32 : NAND4_1 port map( A => L0_31_port, B => L1_31_port, C => 
                           L2_31_port, D => L3_31_port, Y => Y_LOGIC_31_port);
   SHIFTER : BARREL_SHIFTER_N32 port map( CONF => n160, DATA1(31) => DATA1(31),
                           DATA1(30) => DATA1(30), DATA1(29) => DATA1(29), 
                           DATA1(28) => DATA1(28), DATA1(27) => DATA1(27), 
                           DATA1(26) => DATA1(26), DATA1(25) => DATA1(25), 
                           DATA1(24) => DATA1(24), DATA1(23) => DATA1(23), 
                           DATA1(22) => DATA1(22), DATA1(21) => DATA1(21), 
                           DATA1(20) => DATA1(20), DATA1(19) => DATA1(19), 
                           DATA1(18) => DATA1(18), DATA1(17) => DATA1(17), 
                           DATA1(16) => DATA1(16), DATA1(15) => DATA1(15), 
                           DATA1(14) => DATA1(14), DATA1(13) => DATA1(13), 
                           DATA1(12) => DATA1(12), DATA1(11) => DATA1(11), 
                           DATA1(10) => DATA1(10), DATA1(9) => DATA1(9), 
                           DATA1(8) => DATA1(8), DATA1(7) => DATA1(7), DATA1(6)
                           => DATA1(6), DATA1(5) => DATA1(5), DATA1(4) => 
                           DATA1(4), DATA1(3) => DATA1(3), DATA1(2) => DATA1(2)
                           , DATA1(1) => DATA1(1), DATA1(0) => DATA1(0), 
                           DATA2(31) => DATA2(31), DATA2(30) => DATA2(30), 
                           DATA2(29) => DATA2(29), DATA2(28) => DATA2(28), 
                           DATA2(27) => DATA2(27), DATA2(26) => DATA2(26), 
                           DATA2(25) => DATA2(25), DATA2(24) => DATA2(24), 
                           DATA2(23) => DATA2(23), DATA2(22) => DATA2(22), 
                           DATA2(21) => DATA2(21), DATA2(20) => DATA2(20), 
                           DATA2(19) => DATA2(19), DATA2(18) => DATA2(18), 
                           DATA2(17) => DATA2(17), DATA2(16) => DATA2(16), 
                           DATA2(15) => DATA2(15), DATA2(14) => DATA2(14), 
                           DATA2(13) => DATA2(13), DATA2(12) => DATA2(12), 
                           DATA2(11) => DATA2(11), DATA2(10) => DATA2(10), 
                           DATA2(9) => DATA2(9), DATA2(8) => DATA2(8), DATA2(7)
                           => DATA2(7), DATA2(6) => DATA2(6), DATA2(5) => 
                           DATA2(5), DATA2(4) => DATA2(4), DATA2(3) => DATA2(3)
                           , DATA2(2) => DATA2(2), DATA2(1) => DATA2(1), 
                           DATA2(0) => DATA2(0), OUTPUT(31) => 
                           OUT_SHIFTER_31_port, OUTPUT(30) => 
                           OUT_SHIFTER_30_port, OUTPUT(29) => 
                           OUT_SHIFTER_29_port, OUTPUT(28) => 
                           OUT_SHIFTER_28_port, OUTPUT(27) => 
                           OUT_SHIFTER_27_port, OUTPUT(26) => 
                           OUT_SHIFTER_26_port, OUTPUT(25) => 
                           OUT_SHIFTER_25_port, OUTPUT(24) => 
                           OUT_SHIFTER_24_port, OUTPUT(23) => 
                           OUT_SHIFTER_23_port, OUTPUT(22) => 
                           OUT_SHIFTER_22_port, OUTPUT(21) => 
                           OUT_SHIFTER_21_port, OUTPUT(20) => 
                           OUT_SHIFTER_20_port, OUTPUT(19) => 
                           OUT_SHIFTER_19_port, OUTPUT(18) => 
                           OUT_SHIFTER_18_port, OUTPUT(17) => 
                           OUT_SHIFTER_17_port, OUTPUT(16) => 
                           OUT_SHIFTER_16_port, OUTPUT(15) => 
                           OUT_SHIFTER_15_port, OUTPUT(14) => 
                           OUT_SHIFTER_14_port, OUTPUT(13) => 
                           OUT_SHIFTER_13_port, OUTPUT(12) => 
                           OUT_SHIFTER_12_port, OUTPUT(11) => 
                           OUT_SHIFTER_11_port, OUTPUT(10) => 
                           OUT_SHIFTER_10_port, OUTPUT(9) => OUT_SHIFTER_9_port
                           , OUTPUT(8) => OUT_SHIFTER_8_port, OUTPUT(7) => 
                           OUT_SHIFTER_7_port, OUTPUT(6) => OUT_SHIFTER_6_port,
                           OUTPUT(5) => OUT_SHIFTER_5_port, OUTPUT(4) => 
                           OUT_SHIFTER_4_port, OUTPUT(3) => OUT_SHIFTER_3_port,
                           OUTPUT(2) => OUT_SHIFTER_2_port, OUTPUT(1) => 
                           OUT_SHIFTER_1_port, OUTPUT(0) => OUT_SHIFTER_0_port)
                           ;
   r75 : ALU_N32_DW01_addsub_0 port map( A(31) => DATA1(31), A(30) => DATA1(30)
                           , A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , CI => n12, ADD_SUB => U2_U1_Z_0, SUM(31) => N110, 
                           SUM(30) => N109, SUM(29) => N108, SUM(28) => N107, 
                           SUM(27) => N106, SUM(26) => N105, SUM(25) => N104, 
                           SUM(24) => N103, SUM(23) => N102, SUM(22) => N101, 
                           SUM(21) => N100, SUM(20) => N99, SUM(19) => N98, 
                           SUM(18) => N97, SUM(17) => N96, SUM(16) => N95, 
                           SUM(15) => N94, SUM(14) => N93, SUM(13) => N92, 
                           SUM(12) => N91, SUM(11) => N90, SUM(10) => N89, 
                           SUM(9) => N88, SUM(8) => N87, SUM(7) => N86, SUM(6) 
                           => N85, SUM(5) => N84, SUM(4) => N83, SUM(3) => N82,
                           SUM(2) => N81, SUM(1) => N80, SUM(0) => N79, CO => 
                           n_1040);
   r69 : ALU_N32_DW01_cmp6_0 port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , TC => U2_U2_Z_0, LT => n_1041, GT => n_1042, EQ =>
                           n_1043, LE => N111, GE => N112, NE => N113);
   U3 : INV_X4 port map( A => n38, ZN => S_2_port);
   U4 : NAND2_X2 port map( A1 => n38, A2 => n39, ZN => n4);
   U5 : NAND2_X2 port map( A1 => n37, A2 => n46, ZN => n3);
   U6 : NAND2_X2 port map( A1 => n36, A2 => n48, ZN => n2);
   U7 : INV_X2 port map( A => n37, ZN => U2_U1_Z_0);
   U8 : OAI21_X4 port map( B1 => FUNC(3), B2 => n38, A => n39, ZN => S_3_port);
   U9 : INV_X1 port map( A => n1, ZN => OUTALU(31));
   U10 : AOI222_X1 port map( A1 => OUT_SHIFTER_31_port, A2 => n2, B1 => N110, 
                           B2 => n3, C1 => Y_LOGIC_31_port, C2 => n4, ZN => n1)
                           ;
   U11 : INV_X1 port map( A => n5, ZN => OUTALU(26));
   U12 : AOI222_X1 port map( A1 => OUT_SHIFTER_26_port, A2 => n2, B1 => N105, 
                           B2 => n3, C1 => Y_LOGIC_26_port, C2 => n4, ZN => n5)
                           ;
   U13 : INV_X1 port map( A => n6, ZN => OUTALU(27));
   U14 : AOI222_X1 port map( A1 => OUT_SHIFTER_27_port, A2 => n2, B1 => N106, 
                           B2 => n3, C1 => Y_LOGIC_27_port, C2 => n4, ZN => n6)
                           ;
   U15 : INV_X1 port map( A => n7, ZN => OUTALU(24));
   U16 : AOI222_X1 port map( A1 => OUT_SHIFTER_24_port, A2 => n2, B1 => N103, 
                           B2 => n3, C1 => Y_LOGIC_24_port, C2 => n4, ZN => n7)
                           ;
   U17 : INV_X1 port map( A => n8, ZN => OUTALU(25));
   U18 : AOI222_X1 port map( A1 => OUT_SHIFTER_25_port, A2 => n2, B1 => N104, 
                           B2 => n3, C1 => Y_LOGIC_25_port, C2 => n4, ZN => n8)
                           ;
   U19 : INV_X1 port map( A => n9, ZN => OUTALU(30));
   U20 : AOI222_X1 port map( A1 => OUT_SHIFTER_30_port, A2 => n2, B1 => N109, 
                           B2 => n3, C1 => Y_LOGIC_30_port, C2 => n4, ZN => n9)
                           ;
   U21 : INV_X1 port map( A => n10, ZN => OUTALU(28));
   U22 : AOI222_X1 port map( A1 => OUT_SHIFTER_28_port, A2 => n2, B1 => N107, 
                           B2 => n3, C1 => Y_LOGIC_28_port, C2 => n4, ZN => n10
                           );
   U23 : INV_X1 port map( A => n11, ZN => OUTALU(29));
   U24 : AOI222_X1 port map( A1 => OUT_SHIFTER_29_port, A2 => n2, B1 => N108, 
                           B2 => n3, C1 => Y_LOGIC_29_port, C2 => n4, ZN => n11
                           );
   U25 : INV_X1 port map( A => n13, ZN => OUTALU(23));
   U26 : AOI222_X1 port map( A1 => OUT_SHIFTER_23_port, A2 => n2, B1 => N102, 
                           B2 => n3, C1 => Y_LOGIC_23_port, C2 => n4, ZN => n13
                           );
   U27 : INV_X1 port map( A => n14, ZN => OUTALU(10));
   U28 : AOI222_X1 port map( A1 => OUT_SHIFTER_10_port, A2 => n2, B1 => N89, B2
                           => n3, C1 => Y_LOGIC_10_port, C2 => n4, ZN => n14);
   U29 : INV_X1 port map( A => n15, ZN => OUTALU(11));
   U30 : AOI222_X1 port map( A1 => OUT_SHIFTER_11_port, A2 => n2, B1 => N90, B2
                           => n3, C1 => Y_LOGIC_11_port, C2 => n4, ZN => n15);
   U31 : INV_X1 port map( A => n16, ZN => OUTALU(8));
   U32 : AOI222_X1 port map( A1 => OUT_SHIFTER_8_port, A2 => n2, B1 => N87, B2 
                           => n3, C1 => Y_LOGIC_8_port, C2 => n4, ZN => n16);
   U33 : INV_X1 port map( A => n17, ZN => OUTALU(9));
   U34 : AOI222_X1 port map( A1 => OUT_SHIFTER_9_port, A2 => n2, B1 => N88, B2 
                           => n3, C1 => Y_LOGIC_9_port, C2 => n4, ZN => n17);
   U35 : INV_X1 port map( A => n18, ZN => OUTALU(14));
   U36 : AOI222_X1 port map( A1 => OUT_SHIFTER_14_port, A2 => n2, B1 => N93, B2
                           => n3, C1 => Y_LOGIC_14_port, C2 => n4, ZN => n18);
   U37 : INV_X1 port map( A => n19, ZN => OUTALU(15));
   U38 : AOI222_X1 port map( A1 => OUT_SHIFTER_15_port, A2 => n2, B1 => N94, B2
                           => n3, C1 => Y_LOGIC_15_port, C2 => n4, ZN => n19);
   U39 : INV_X1 port map( A => n20, ZN => OUTALU(12));
   U40 : AOI222_X1 port map( A1 => OUT_SHIFTER_12_port, A2 => n2, B1 => N91, B2
                           => n3, C1 => Y_LOGIC_12_port, C2 => n4, ZN => n20);
   U41 : INV_X1 port map( A => n21, ZN => OUTALU(13));
   U42 : AOI222_X1 port map( A1 => OUT_SHIFTER_13_port, A2 => n2, B1 => N92, B2
                           => n3, C1 => Y_LOGIC_13_port, C2 => n4, ZN => n21);
   U43 : INV_X1 port map( A => n22, ZN => OUTALU(7));
   U44 : AOI222_X1 port map( A1 => OUT_SHIFTER_7_port, A2 => n2, B1 => N86, B2 
                           => n3, C1 => Y_LOGIC_7_port, C2 => n4, ZN => n22);
   U45 : INV_X1 port map( A => n23, ZN => OUTALU(18));
   U46 : AOI222_X1 port map( A1 => OUT_SHIFTER_18_port, A2 => n2, B1 => N97, B2
                           => n3, C1 => Y_LOGIC_18_port, C2 => n4, ZN => n23);
   U47 : INV_X1 port map( A => n24, ZN => OUTALU(19));
   U48 : AOI222_X1 port map( A1 => OUT_SHIFTER_19_port, A2 => n2, B1 => N98, B2
                           => n3, C1 => Y_LOGIC_19_port, C2 => n4, ZN => n24);
   U49 : INV_X1 port map( A => n25, ZN => OUTALU(16));
   U50 : AOI222_X1 port map( A1 => OUT_SHIFTER_16_port, A2 => n2, B1 => N95, B2
                           => n3, C1 => Y_LOGIC_16_port, C2 => n4, ZN => n25);
   U51 : INV_X1 port map( A => n26, ZN => OUTALU(17));
   U52 : AOI222_X1 port map( A1 => OUT_SHIFTER_17_port, A2 => n2, B1 => N96, B2
                           => n3, C1 => Y_LOGIC_17_port, C2 => n4, ZN => n26);
   U53 : INV_X1 port map( A => n27, ZN => OUTALU(22));
   U54 : AOI222_X1 port map( A1 => OUT_SHIFTER_22_port, A2 => n2, B1 => N101, 
                           B2 => n3, C1 => Y_LOGIC_22_port, C2 => n4, ZN => n27
                           );
   U55 : INV_X1 port map( A => n28, ZN => OUTALU(20));
   U56 : AOI222_X1 port map( A1 => OUT_SHIFTER_20_port, A2 => n2, B1 => N99, B2
                           => n3, C1 => Y_LOGIC_20_port, C2 => n4, ZN => n28);
   U57 : INV_X1 port map( A => n29, ZN => OUTALU(21));
   U58 : AOI222_X1 port map( A1 => OUT_SHIFTER_21_port, A2 => n2, B1 => N100, 
                           B2 => n3, C1 => Y_LOGIC_21_port, C2 => n4, ZN => n29
                           );
   U59 : INV_X1 port map( A => n30, ZN => OUTALU(2));
   U60 : AOI222_X1 port map( A1 => OUT_SHIFTER_2_port, A2 => n2, B1 => N81, B2 
                           => n3, C1 => Y_LOGIC_2_port, C2 => n4, ZN => n30);
   U61 : INV_X1 port map( A => n31, ZN => OUTALU(3));
   U62 : AOI222_X1 port map( A1 => OUT_SHIFTER_3_port, A2 => n2, B1 => N82, B2 
                           => n3, C1 => Y_LOGIC_3_port, C2 => n4, ZN => n31);
   U63 : INV_X1 port map( A => n32, ZN => OUTALU(1));
   U64 : AOI222_X1 port map( A1 => OUT_SHIFTER_1_port, A2 => n2, B1 => N80, B2 
                           => n3, C1 => Y_LOGIC_1_port, C2 => n4, ZN => n32);
   U65 : INV_X1 port map( A => n33, ZN => OUTALU(6));
   U66 : AOI222_X1 port map( A1 => OUT_SHIFTER_6_port, A2 => n2, B1 => N85, B2 
                           => n3, C1 => Y_LOGIC_6_port, C2 => n4, ZN => n33);
   U67 : INV_X1 port map( A => n34, ZN => OUTALU(4));
   U68 : AOI222_X1 port map( A1 => OUT_SHIFTER_4_port, A2 => n2, B1 => N83, B2 
                           => n3, C1 => Y_LOGIC_4_port, C2 => n4, ZN => n34);
   U69 : INV_X1 port map( A => n35, ZN => OUTALU(5));
   U70 : AOI222_X1 port map( A1 => OUT_SHIFTER_5_port, A2 => n2, B1 => N84, B2 
                           => n3, C1 => Y_LOGIC_5_port, C2 => n4, ZN => n35);
   U71 : INV_X1 port map( A => DATA1(31), ZN => n84_port);
   U72 : INV_X1 port map( A => DATA1(30), ZN => n85_port);
   U73 : INV_X1 port map( A => DATA1(29), ZN => n86_port);
   U74 : INV_X1 port map( A => DATA1(28), ZN => n87_port);
   U75 : INV_X1 port map( A => DATA1(27), ZN => n88_port);
   U76 : INV_X1 port map( A => DATA1(26), ZN => n89_port);
   U77 : INV_X1 port map( A => DATA1(25), ZN => n90_port);
   U78 : INV_X1 port map( A => DATA1(24), ZN => n91_port);
   U79 : INV_X1 port map( A => DATA1(23), ZN => n92_port);
   U80 : INV_X1 port map( A => DATA1(22), ZN => n93_port);
   U81 : INV_X1 port map( A => DATA1(21), ZN => n94_port);
   U82 : INV_X1 port map( A => DATA1(20), ZN => n95_port);
   U83 : INV_X1 port map( A => DATA1(19), ZN => n96_port);
   U84 : INV_X1 port map( A => DATA1(18), ZN => n97_port);
   U85 : INV_X1 port map( A => DATA1(17), ZN => n98_port);
   U86 : INV_X1 port map( A => DATA1(16), ZN => n99_port);
   U87 : INV_X1 port map( A => DATA1(15), ZN => n100_port);
   U88 : INV_X1 port map( A => DATA1(14), ZN => n101_port);
   U89 : INV_X1 port map( A => DATA1(13), ZN => n102_port);
   U90 : INV_X1 port map( A => DATA1(12), ZN => n103_port);
   U91 : INV_X1 port map( A => DATA1(11), ZN => n104_port);
   U92 : INV_X1 port map( A => DATA1(10), ZN => n105_port);
   U93 : INV_X1 port map( A => DATA1(9), ZN => n106_port);
   U94 : INV_X1 port map( A => DATA1(8), ZN => n107_port);
   U95 : INV_X1 port map( A => DATA1(7), ZN => n108_port);
   U96 : INV_X1 port map( A => DATA1(6), ZN => n109_port);
   U97 : INV_X1 port map( A => DATA1(5), ZN => n110_port);
   U98 : INV_X1 port map( A => DATA1(4), ZN => n111_port);
   U99 : INV_X1 port map( A => DATA1(3), ZN => n112_port);
   U100 : INV_X1 port map( A => DATA1(2), ZN => n113_port);
   U101 : INV_X1 port map( A => DATA1(1), ZN => n114);
   U102 : INV_X1 port map( A => DATA1(0), ZN => n115);
   U103 : INV_X1 port map( A => DATA2(31), ZN => n116);
   U104 : INV_X1 port map( A => DATA2(30), ZN => n117);
   U105 : INV_X1 port map( A => DATA2(29), ZN => n118);
   U106 : INV_X1 port map( A => DATA2(28), ZN => n119);
   U107 : INV_X1 port map( A => DATA2(27), ZN => n120);
   U108 : INV_X1 port map( A => DATA2(26), ZN => n121);
   U109 : INV_X1 port map( A => DATA2(25), ZN => n122);
   U110 : INV_X1 port map( A => DATA2(24), ZN => n123);
   U111 : INV_X1 port map( A => DATA2(23), ZN => n124);
   U112 : INV_X1 port map( A => DATA2(22), ZN => n125);
   U113 : INV_X1 port map( A => DATA2(21), ZN => n126);
   U114 : INV_X1 port map( A => DATA2(20), ZN => n127);
   U115 : INV_X1 port map( A => DATA2(19), ZN => n128);
   U116 : INV_X1 port map( A => DATA2(18), ZN => n129);
   U117 : INV_X1 port map( A => DATA2(17), ZN => n130);
   U118 : INV_X1 port map( A => DATA2(16), ZN => n131);
   U119 : INV_X1 port map( A => DATA2(15), ZN => n132);
   U120 : INV_X1 port map( A => DATA2(14), ZN => n133);
   U121 : INV_X1 port map( A => DATA2(13), ZN => n134);
   U122 : INV_X1 port map( A => DATA2(12), ZN => n135);
   U123 : INV_X1 port map( A => DATA2(11), ZN => n136);
   U124 : INV_X1 port map( A => DATA2(10), ZN => n137);
   U125 : INV_X1 port map( A => DATA2(9), ZN => n138);
   U126 : INV_X1 port map( A => DATA2(8), ZN => n139);
   U127 : INV_X1 port map( A => DATA2(7), ZN => n140);
   U128 : INV_X1 port map( A => DATA2(6), ZN => n141);
   U129 : INV_X1 port map( A => DATA2(5), ZN => n142);
   U130 : INV_X1 port map( A => DATA2(4), ZN => n143);
   U131 : INV_X1 port map( A => DATA2(3), ZN => n144);
   U132 : INV_X1 port map( A => DATA2(2), ZN => n145);
   U133 : INV_X1 port map( A => DATA2(1), ZN => n146);
   U134 : INV_X1 port map( A => DATA2(0), ZN => n147);
   U135 : INV_X1 port map( A => n36, ZN => n160);
   U136 : NAND3_X1 port map( A1 => n40, A2 => n41, A3 => n42, ZN => OUTALU(0));
   U137 : AOI22_X1 port map( A1 => N79, A2 => n3, B1 => Y_LOGIC_0_port, B2 => 
                           n4, ZN => n42);
   U138 : NAND3_X1 port map( A1 => FUNC(3), A2 => n43, A3 => FUNC(2), ZN => n39
                           );
   U139 : NAND3_X1 port map( A1 => n44, A2 => n45, A3 => FUNC(1), ZN => n38);
   U140 : NAND3_X1 port map( A1 => n43, A2 => n44, A3 => FUNC(3), ZN => n46);
   U141 : NAND3_X1 port map( A1 => n43, A2 => n47, A3 => FUNC(2), ZN => n37);
   U142 : NOR2_X1 port map( A1 => FUNC(1), A2 => FUNC(0), ZN => n43);
   U143 : NAND2_X1 port map( A1 => OUT_SHIFTER_0_port, A2 => n2, ZN => n41);
   U144 : NAND3_X1 port map( A1 => FUNC(2), A2 => n47, A3 => n49, ZN => n48);
   U145 : INV_X1 port map( A => FUNC(3), ZN => n47);
   U146 : NAND3_X1 port map( A1 => FUNC(3), A2 => n44, A3 => n49, ZN => n36);
   U147 : MUX2_X1 port map( A => n50, B => n51, S => FUNC(3), Z => n40);
   U148 : NAND2_X1 port map( A1 => N112, A2 => U2_U2_Z_0, ZN => n51);
   U149 : AOI22_X1 port map( A1 => n52, A2 => N113, B1 => N111, B2 => U2_U2_Z_0
                           , ZN => n50);
   U150 : AND3_X1 port map( A1 => FUNC(2), A2 => n45, A3 => FUNC(1), ZN => 
                           U2_U2_Z_0);
   U151 : AND2_X1 port map( A1 => n44, A2 => n49, ZN => n52);
   U152 : NOR2_X1 port map( A1 => n45, A2 => FUNC(1), ZN => n49);
   U153 : INV_X1 port map( A => FUNC(0), ZN => n45);
   U154 : INV_X1 port map( A => FUNC(2), ZN => n44);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26 is

   port( NOT_EXT_IMM : in std_logic_vector (25 downto 0);  SIGNED_IMM, IS_JUMP 
         : in std_logic;  EXT_IMM : out std_logic_vector (31 downto 0));

end EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26;

architecture SYN_BEHAVIOR of EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal EXT_IMM_31_port, EXT_IMM_25_port, EXT_IMM_24_port, EXT_IMM_23_port, 
      EXT_IMM_22_port, EXT_IMM_21_port, EXT_IMM_20_port, EXT_IMM_19_port, 
      EXT_IMM_18_port, EXT_IMM_17_port, EXT_IMM_16_port, n1, n2, n3, n4, n5, n6
      , n7, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   EXT_IMM <= ( EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, 
      EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_31_port, EXT_IMM_25_port, 
      EXT_IMM_24_port, EXT_IMM_23_port, EXT_IMM_22_port, EXT_IMM_21_port, 
      EXT_IMM_20_port, EXT_IMM_19_port, EXT_IMM_18_port, EXT_IMM_17_port, 
      EXT_IMM_16_port, NOT_EXT_IMM(15), NOT_EXT_IMM(14), NOT_EXT_IMM(13), 
      NOT_EXT_IMM(12), NOT_EXT_IMM(11), NOT_EXT_IMM(10), NOT_EXT_IMM(9), 
      NOT_EXT_IMM(8), NOT_EXT_IMM(7), NOT_EXT_IMM(6), NOT_EXT_IMM(5), 
      NOT_EXT_IMM(4), NOT_EXT_IMM(3), NOT_EXT_IMM(2), NOT_EXT_IMM(1), 
      NOT_EXT_IMM(0) );
   
   U2 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => EXT_IMM_31_port);
   U3 : NAND3_X1 port map( A1 => NOT_EXT_IMM(25), A2 => IS_JUMP, A3 => 
                           SIGNED_IMM, ZN => n2);
   U4 : OAI21_X1 port map( B1 => n3, B2 => n4, A => n1, ZN => EXT_IMM_25_port);
   U5 : INV_X1 port map( A => NOT_EXT_IMM(25), ZN => n4);
   U6 : NAND2_X1 port map( A1 => n1, A2 => n5, ZN => EXT_IMM_24_port);
   U7 : NAND2_X1 port map( A1 => NOT_EXT_IMM(24), A2 => IS_JUMP, ZN => n5);
   U8 : NAND2_X1 port map( A1 => n1, A2 => n6, ZN => EXT_IMM_23_port);
   U9 : NAND2_X1 port map( A1 => NOT_EXT_IMM(23), A2 => IS_JUMP, ZN => n6);
   U10 : NAND2_X1 port map( A1 => n1, A2 => n7, ZN => EXT_IMM_22_port);
   U11 : NAND2_X1 port map( A1 => NOT_EXT_IMM(22), A2 => IS_JUMP, ZN => n7);
   U12 : NAND2_X1 port map( A1 => n1, A2 => n8, ZN => EXT_IMM_21_port);
   U13 : NAND2_X1 port map( A1 => NOT_EXT_IMM(21), A2 => IS_JUMP, ZN => n8);
   U14 : NAND2_X1 port map( A1 => n1, A2 => n9, ZN => EXT_IMM_20_port);
   U15 : NAND2_X1 port map( A1 => NOT_EXT_IMM(20), A2 => IS_JUMP, ZN => n9);
   U16 : NAND2_X1 port map( A1 => n1, A2 => n10, ZN => EXT_IMM_19_port);
   U17 : NAND2_X1 port map( A1 => NOT_EXT_IMM(19), A2 => IS_JUMP, ZN => n10);
   U18 : NAND2_X1 port map( A1 => n1, A2 => n11, ZN => EXT_IMM_18_port);
   U19 : NAND2_X1 port map( A1 => NOT_EXT_IMM(18), A2 => IS_JUMP, ZN => n11);
   U20 : NAND2_X1 port map( A1 => n1, A2 => n12, ZN => EXT_IMM_17_port);
   U21 : NAND2_X1 port map( A1 => NOT_EXT_IMM(17), A2 => IS_JUMP, ZN => n12);
   U22 : NAND2_X1 port map( A1 => n1, A2 => n13, ZN => EXT_IMM_16_port);
   U23 : NAND2_X1 port map( A1 => NOT_EXT_IMM(16), A2 => IS_JUMP, ZN => n13);
   U24 : NAND3_X1 port map( A1 => SIGNED_IMM, A2 => n3, A3 => NOT_EXT_IMM(15), 
                           ZN => n1);
   U25 : INV_X1 port map( A => IS_JUMP, ZN => n3);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REGISTER_FILE_NBIT32_NREG32 is

   port( CLK, RST, EN, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 :
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0));

end REGISTER_FILE_NBIT32_NREG32;

architecture SYN_BEHAVIOR of REGISTER_FILE_NBIT32_NREG32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n833, n834, n835, n836, n837, n838, n839, 
      n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, 
      n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
      n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
      n888, n889, n890, n891, n892, n893, n894, n895, n896, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n2527, n2528, n2529, n2530, n2531, 
      n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, 
      n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, 
      n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, 
      n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, 
      n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, 
      n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
      n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, 
      n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, 
      n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, 
      n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
      n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, 
      n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, 
      n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, 
      n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, 
      n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, 
      n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, 
      n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, 
      n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, 
      n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, 
      n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, 
      n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, 
      n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, 
      n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, 
      n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, 
      n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, 
      n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, 
      n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, 
      n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, 
      n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, 
      n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, 
      n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, 
      n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, 
      n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, 
      n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, 
      n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, 
      n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
      n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
      n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, 
      n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
      n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, 
      n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, 
      n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, 
      n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, 
      n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, 
      n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
      n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, 
      n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
      n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, 
      n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, 
      n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, 
      n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, 
      n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, 
      n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, 
      n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, 
      n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
      n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
      n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
      n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, 
      n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
      n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
      n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, 
      n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, 
      n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, 
      n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, 
      n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, 
      n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, 
      n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
      n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
      n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, 
      n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, 
      n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, 
      n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, 
      n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, 
      n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, 
      n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
      n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, 
      n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, 
      n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, 
      n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, 
      n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, 
      n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, 
      n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, 
      n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, 
      n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, 
      n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, 
      n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, 
      n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, 
      n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, 
      n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, 
      n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, 
      n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, 
      n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, 
      n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, 
      n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, 
      n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, 
      n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, 
      n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, 
      n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, 
      n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, 
      n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, 
      n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, 
      n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, 
      n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, 
      n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, 
      n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, 
      n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, 
      n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, 
      n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, 
      n3612, n3613, n3614, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, 
      n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
      n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n507, n508, n509, n510, n511, n512, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, 
      n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
      n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, 
      n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, 
      n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, 
      n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, 
      n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, 
      n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, 
      n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, 
      n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, 
      n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, 
      n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, 
      n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, 
      n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, 
      n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, 
      n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, 
      n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, 
      n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, 
      n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, 
      n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, 
      n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, 
      n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, 
      n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, 
      n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, 
      n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, 
      n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, 
      n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, 
      n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, 
      n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, 
      n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, 
      n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
      n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, 
      n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, 
      n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, 
      n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, 
      n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, 
      n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, 
      n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, 
      n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, 
      n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, 
      n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, 
      n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, 
      n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, 
      n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, 
      n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, 
      n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, 
      n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, 
      n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, 
      n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, 
      n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, 
      n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, 
      n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, 
      n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, 
      n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
      n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, 
      n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, 
      n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, 
      n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, 
      n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, 
      n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, 
      n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
      n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, 
      n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, 
      n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, 
      n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, 
      n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, 
      n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, 
      n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, 
      n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, 
      n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, 
      n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, 
      n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, 
      n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, 
      n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, 
      n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, 
      n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, 
      n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, 
      n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, 
      n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, 
      n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, 
      n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, 
      n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, 
      n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, 
      n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, 
      n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, 
      n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
      n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, 
      n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, 
      n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, 
      n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, 
      n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, 
      n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, 
      n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, 
      n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, 
      n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, 
      n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, 
      n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, 
      n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, 
      n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, 
      n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, 
      n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, 
      n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, 
      n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, 
      n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, 
      n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, 
      n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, 
      n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
      n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, 
      n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, 
      n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, 
      n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, 
      n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, 
      n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, 
      n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, 
      n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, 
      n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, 
      n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, 
      n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, 
      n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, 
      n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, 
      n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, 
      n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, 
      n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, 
      n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, 
      n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, 
      n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, 
      n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, 
      n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, 
      n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, 
      n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, 
      n2524, n2525, n2526, n3615, n3616, n3617, n3618, n3619, n3620, n3621, 
      n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, 
      n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, 
      n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, 
      n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, 
      n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, 
      n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, 
      n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, 
      n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, 
      n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, 
      n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, 
      n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, 
      n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, 
      n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, 
      n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, 
      n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, 
      n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, 
      n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, 
      n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, 
      n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, 
      n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, 
      n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, 
      n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, 
      n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, 
      n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, 
      n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, 
      n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, 
      n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, 
      n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, 
      n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, 
      n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, 
      n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, 
      n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, 
      n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, 
      n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, 
      n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, 
      n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, 
      n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, 
      n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, 
      n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, 
      n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, 
      n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, 
      n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, 
      n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, 
      n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, 
      n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, 
      n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, 
      n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, 
      n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, 
      n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, 
      n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, 
      n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, 
      n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, 
      n4142, n4143, n4144, n4145, n4146, n4147, n4148, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n3614, CK => CLK, Q => n130,
                           QN => n_1044);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => n132,
                           QN => n_1045);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => n134,
                           QN => n_1046);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => n136,
                           QN => n_1047);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => n138,
                           QN => n_1048);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => n140,
                           QN => n_1049);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => n142,
                           QN => n_1050);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => n144,
                           QN => n_1051);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => n146,
                           QN => n_1052);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => n148,
                           QN => n_1053);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => n150,
                           QN => n_1054);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => n152,
                           QN => n_1055);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => n154,
                           QN => n_1056);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => n156,
                           QN => n_1057);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => n158,
                           QN => n_1058);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => n160,
                           QN => n_1059);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => n162,
                           QN => n_1060);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => n164,
                           QN => n_1061);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => n166,
                           QN => n_1062);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => n168,
                           QN => n_1063);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => n170,
                           QN => n_1064);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => n172,
                           QN => n_1065);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => n174, 
                           QN => n_1066);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => n176, 
                           QN => n_1067);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => n178, 
                           QN => n_1068);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => n180, 
                           QN => n_1069);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => n182, 
                           QN => n_1070);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => n184, 
                           QN => n_1071);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => n186, 
                           QN => n_1072);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => n188, 
                           QN => n_1073);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => n190, 
                           QN => n_1074);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => n192, 
                           QN => n_1075);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => n2, 
                           QN => n_1076);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => n4, 
                           QN => n_1077);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => n6, 
                           QN => n_1078);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => n8, 
                           QN => n_1079);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => n10, 
                           QN => n_1080);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => n12, 
                           QN => n_1081);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => n14, 
                           QN => n_1082);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => n16, 
                           QN => n_1083);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => n18, 
                           QN => n_1084);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => n20, 
                           QN => n_1085);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => n22, 
                           QN => n_1086);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => n24, 
                           QN => n_1087);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => n26, 
                           QN => n_1088);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => n28, 
                           QN => n_1089);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => n30, 
                           QN => n_1090);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => n32, 
                           QN => n_1091);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => n34, 
                           QN => n_1092);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => n36, 
                           QN => n_1093);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => n38, 
                           QN => n_1094);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => n40, 
                           QN => n_1095);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => n42, 
                           QN => n_1096);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => n44, 
                           QN => n_1097);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => n46, 
                           QN => n_1098);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => n48, 
                           QN => n_1099);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => n50, 
                           QN => n_1100);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => n52, 
                           QN => n_1101);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => n54, 
                           QN => n_1102);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => n56, 
                           QN => n_1103);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => n58, 
                           QN => n_1104);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => n60, 
                           QN => n_1105);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => n62, 
                           QN => n_1106);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => n64, 
                           QN => n_1107);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => n4148
                           , QN => n66);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => n4147
                           , QN => n68);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => n4146
                           , QN => n70);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => n4145
                           , QN => n72);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => n4144
                           , QN => n74);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => n4143
                           , QN => n76);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => n4142
                           , QN => n78);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => n4141
                           , QN => n80);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => n4140
                           , QN => n82);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => n4139
                           , QN => n84);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => n4138
                           , QN => n86);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => n4137
                           , QN => n88);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => n4136
                           , QN => n90);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => n4135
                           , QN => n92);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => n4134
                           , QN => n94);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => n4133
                           , QN => n96);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => n4132
                           , QN => n98);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => n4131
                           , QN => n100);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => n4130
                           , QN => n102);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => n4129
                           , QN => n104);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => n4128
                           , QN => n106);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => n4127
                           , QN => n108);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => n4126,
                           QN => n110);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => n4125,
                           QN => n112);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n3526, CK => CLK, Q => n4124,
                           QN => n114);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => n4123,
                           QN => n116);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => n4122,
                           QN => n118);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => n4121,
                           QN => n120);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => n4120,
                           QN => n122);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => n4119,
                           QN => n124);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => n4118,
                           QN => n126);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => n4117,
                           QN => n128);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => n4116
                           , QN => n194);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => n4115
                           , QN => n196);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => n4114
                           , QN => n198);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => n4113
                           , QN => n200);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => n4112
                           , QN => n202);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => n4111
                           , QN => n204);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => n4110
                           , QN => n206);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => n4109
                           , QN => n208);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => n4108
                           , QN => n210);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => n4107
                           , QN => n212);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => n4106
                           , QN => n214);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => n4105
                           , QN => n216);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => n4104
                           , QN => n218);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => n4103
                           , QN => n220);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => n4102
                           , QN => n222);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => n4101
                           , QN => n224);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => n4100
                           , QN => n226);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => n4099
                           , QN => n228);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => n4098
                           , QN => n230);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => n4097
                           , QN => n232);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => n4096
                           , QN => n234);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => n4095
                           , QN => n236);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => n4094,
                           QN => n238);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => n4093,
                           QN => n240);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => n4092,
                           QN => n242);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => n4091,
                           QN => n244);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => n4090,
                           QN => n246);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => n4089,
                           QN => n248);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => n4088,
                           QN => n250);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => n4087,
                           QN => n252);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => n4086,
                           QN => n254);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => n4085,
                           QN => n256);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => n129,
                           QN => n_1108);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => n131,
                           QN => n_1109);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => n133,
                           QN => n_1110);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => n135,
                           QN => n_1111);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => n137,
                           QN => n_1112);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => n139,
                           QN => n_1113);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => n141,
                           QN => n_1114);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => n143,
                           QN => n_1115);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => n145,
                           QN => n_1116);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => n147,
                           QN => n_1117);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => n149,
                           QN => n_1118);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => n151,
                           QN => n_1119);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => n153,
                           QN => n_1120);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => n155,
                           QN => n_1121);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n3472, CK => CLK, Q => n157,
                           QN => n_1122);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => n159,
                           QN => n_1123);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => n161,
                           QN => n_1124);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => n163,
                           QN => n_1125);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => n165,
                           QN => n_1126);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => n167,
                           QN => n_1127);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => n169,
                           QN => n_1128);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => n171,
                           QN => n_1129);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => n173, 
                           QN => n_1130);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => n175, 
                           QN => n_1131);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => n177, 
                           QN => n_1132);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => n179, 
                           QN => n_1133);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => n181, 
                           QN => n_1134);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => n183, 
                           QN => n_1135);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => n185, 
                           QN => n_1136);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => n187, 
                           QN => n_1137);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => n189, 
                           QN => n_1138);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => n191, 
                           QN => n_1139);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => n1, 
                           QN => n_1140);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => n3, 
                           QN => n_1141);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => n5, 
                           QN => n_1142);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => n7, 
                           QN => n_1143);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => n9, 
                           QN => n_1144);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => n11, 
                           QN => n_1145);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => n13, 
                           QN => n_1146);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => n15, 
                           QN => n_1147);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => n17, 
                           QN => n_1148);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => n19, 
                           QN => n_1149);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => n21, 
                           QN => n_1150);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => n23, 
                           QN => n_1151);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => n25, 
                           QN => n_1152);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => n27, 
                           QN => n_1153);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => n29, 
                           QN => n_1154);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => n31, 
                           QN => n_1155);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => n33, 
                           QN => n_1156);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => n35, 
                           QN => n_1157);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => n37, 
                           QN => n_1158);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => n39, 
                           QN => n_1159);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => n41, 
                           QN => n_1160);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => n43, 
                           QN => n_1161);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => n45, 
                           QN => n_1162);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => n47, 
                           QN => n_1163);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => n49, 
                           QN => n_1164);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => n51, 
                           QN => n_1165);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => n53, 
                           QN => n_1166);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => n55, 
                           QN => n_1167);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => n57, 
                           QN => n_1168);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => n59, 
                           QN => n_1169);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => n61, 
                           QN => n_1170);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => n63, 
                           QN => n_1171);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => n4084
                           , QN => n65);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => n4083
                           , QN => n67);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => n4082
                           , QN => n69);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => n4081
                           , QN => n71);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => n4080
                           , QN => n73);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => n4079
                           , QN => n75);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => n4078
                           , QN => n77);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => n4077
                           , QN => n79);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => n4076
                           , QN => n81);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => n4075
                           , QN => n83);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => n4074
                           , QN => n85);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => n4073
                           , QN => n87);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => n4072
                           , QN => n89);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => n4071
                           , QN => n91);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => n4070
                           , QN => n93);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => n4069
                           , QN => n95);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => n4068
                           , QN => n97);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => n4067
                           , QN => n99);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => n4066
                           , QN => n101);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => n4065
                           , QN => n103);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => n4064
                           , QN => n105);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => n4063
                           , QN => n107);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => n4062,
                           QN => n109);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => n4061,
                           QN => n111);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => n4060,
                           QN => n113);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => n4059,
                           QN => n115);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => n4058,
                           QN => n117);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => n4057,
                           QN => n119);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => n4056,
                           QN => n121);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => n4055,
                           QN => n123);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => n4054,
                           QN => n125);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => n4053,
                           QN => n127);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => n4052
                           , QN => n193);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => n4051
                           , QN => n195);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => n4050
                           , QN => n197);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => n4049
                           , QN => n199);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => n4048
                           , QN => n201);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => n4047
                           , QN => n203);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => n4046
                           , QN => n205);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => n4045
                           , QN => n207);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => n4044
                           , QN => n209);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => n4043
                           , QN => n211);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => n4042
                           , QN => n213);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => n4041
                           , QN => n215);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => n4040
                           , QN => n217);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => n4039
                           , QN => n219);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => n4038
                           , QN => n221);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => n4037
                           , QN => n223);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => n4036
                           , QN => n225);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => n4035
                           , QN => n227);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => n4034
                           , QN => n229);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => n4033
                           , QN => n231);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => n4032
                           , QN => n233);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => n4031
                           , QN => n235);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => n4030,
                           QN => n237);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => n4029,
                           QN => n239);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => n4028,
                           QN => n241);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => n4027,
                           QN => n243);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => n4026,
                           QN => n245);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => n4025,
                           QN => n247);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => n4024,
                           QN => n249);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => n4023,
                           QN => n251);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => n4022,
                           QN => n253);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => n4021,
                           QN => n255);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => n705,
                           QN => n257);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => n706,
                           QN => n258);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => n707,
                           QN => n259);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => n708,
                           QN => n260);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => n709,
                           QN => n261);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => n710,
                           QN => n262);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => n711,
                           QN => n263);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => n712,
                           QN => n264);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => n713,
                           QN => n265);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => n714,
                           QN => n266);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => n715,
                           QN => n267);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => n716,
                           QN => n268);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => n717,
                           QN => n269);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => n718,
                           QN => n270);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => n719,
                           QN => n271);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => n720,
                           QN => n272);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => n721,
                           QN => n273);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => n722,
                           QN => n274);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => n723,
                           QN => n275);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => n724,
                           QN => n276);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => n725,
                           QN => n277);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => n726,
                           QN => n278);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => n727, 
                           QN => n279);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => n728, 
                           QN => n280);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => n729, 
                           QN => n281);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => n730, 
                           QN => n282);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => n731, 
                           QN => n283);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => n732, 
                           QN => n284);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => n733, 
                           QN => n285);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => n734, 
                           QN => n286);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => n735, 
                           QN => n287);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => n736, 
                           QN => n288);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3326, CK => CLK, Q => n321,
                           QN => n289);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => n322,
                           QN => n290);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => n323,
                           QN => n291);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => n324,
                           QN => n292);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => n325,
                           QN => n293);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => n326,
                           QN => n294);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => n327,
                           QN => n295);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => n328,
                           QN => n296);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => n329,
                           QN => n297);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => n330,
                           QN => n298);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => n331,
                           QN => n299);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => n332,
                           QN => n300);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => n333,
                           QN => n301);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => n334,
                           QN => n302);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => n335,
                           QN => n303);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => n336,
                           QN => n304);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => n337,
                           QN => n305);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => n338,
                           QN => n306);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => n339,
                           QN => n307);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => n340,
                           QN => n308);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => n341,
                           QN => n309);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => n342,
                           QN => n310);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => n343, 
                           QN => n311);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => n344, 
                           QN => n312);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => n345, 
                           QN => n313);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => n346, 
                           QN => n314);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => n347, 
                           QN => n315);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => n348, 
                           QN => n316);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => n349, 
                           QN => n317);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => n350, 
                           QN => n318);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => n351, 
                           QN => n319);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => n352, 
                           QN => n320);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => 
                           n4020, QN => n_1172);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => 
                           n4019, QN => n_1173);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => 
                           n4018, QN => n_1174);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => 
                           n4017, QN => n_1175);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => 
                           n4016, QN => n_1176);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3289, CK => CLK, Q => 
                           n4015, QN => n_1177);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => 
                           n4014, QN => n_1178);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => 
                           n4013, QN => n_1179);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => 
                           n4012, QN => n_1180);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => 
                           n4011, QN => n_1181);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => 
                           n4010, QN => n_1182);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => 
                           n4009, QN => n_1183);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => 
                           n4008, QN => n_1184);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => 
                           n4007, QN => n_1185);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => 
                           n4006, QN => n_1186);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => 
                           n4005, QN => n_1187);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => 
                           n4004, QN => n_1188);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => 
                           n4003, QN => n_1189);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => 
                           n4002, QN => n_1190);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => 
                           n4001, QN => n_1191);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3274, CK => CLK, Q => 
                           n4000, QN => n_1192);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3273, CK => CLK, Q => 
                           n3999, QN => n_1193);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3272, CK => CLK, Q => n3998
                           , QN => n_1194);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3271, CK => CLK, Q => n3997
                           , QN => n_1195);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3270, CK => CLK, Q => n3996
                           , QN => n_1196);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3269, CK => CLK, Q => n3995
                           , QN => n_1197);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3268, CK => CLK, Q => n3994
                           , QN => n_1198);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3267, CK => CLK, Q => n3993
                           , QN => n_1199);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3266, CK => CLK, Q => n3992
                           , QN => n_1200);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3265, CK => CLK, Q => n3991
                           , QN => n_1201);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3264, CK => CLK, Q => n3990
                           , QN => n_1202);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3263, CK => CLK, Q => n3989
                           , QN => n_1203);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3262, CK => CLK, Q => 
                           n3988, QN => n_1204);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => 
                           n3987, QN => n_1205);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => 
                           n3986, QN => n_1206);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => 
                           n3985, QN => n_1207);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => 
                           n3984, QN => n_1208);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => 
                           n3983, QN => n_1209);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => 
                           n3982, QN => n_1210);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => 
                           n3981, QN => n_1211);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => 
                           n3980, QN => n_1212);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => 
                           n3979, QN => n_1213);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => 
                           n3978, QN => n_1214);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => 
                           n3977, QN => n_1215);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => 
                           n3976, QN => n_1216);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => 
                           n3975, QN => n_1217);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => 
                           n3974, QN => n_1218);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => 
                           n3973, QN => n_1219);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => 
                           n3972, QN => n_1220);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => 
                           n3971, QN => n_1221);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => 
                           n3970, QN => n_1222);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => 
                           n3969, QN => n_1223);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => 
                           n3968, QN => n_1224);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => 
                           n3967, QN => n_1225);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => n3966
                           , QN => n_1226);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => n3965
                           , QN => n_1227);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => n3964
                           , QN => n_1228);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => n3963
                           , QN => n_1229);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => n3962
                           , QN => n_1230);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => n3961
                           , QN => n_1231);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => n3960
                           , QN => n_1232);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => n3959
                           , QN => n_1233);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => n3958
                           , QN => n_1234);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => n3957
                           , QN => n_1235);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => n737
                           , QN => n385);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => n738
                           , QN => n386);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => n739
                           , QN => n387);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => n740
                           , QN => n388);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => n741
                           , QN => n389);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => n742
                           , QN => n390);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => n743
                           , QN => n391);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => n744
                           , QN => n392);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => n745
                           , QN => n393);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => n746
                           , QN => n394);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => n747
                           , QN => n395);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => n748
                           , QN => n396);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => n749
                           , QN => n397);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => n750
                           , QN => n398);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => n751
                           , QN => n399);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => n752
                           , QN => n400);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => n753
                           , QN => n401);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => n754
                           , QN => n402);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => n755
                           , QN => n403);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => n756
                           , QN => n404);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => n757
                           , QN => n405);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => n758
                           , QN => n406);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3208, CK => CLK, Q => n759,
                           QN => n407);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => n760,
                           QN => n408);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => n761,
                           QN => n409);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => n762,
                           QN => n410);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => n763,
                           QN => n411);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => n764,
                           QN => n412);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => n765,
                           QN => n413);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => n766,
                           QN => n414);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => n767,
                           QN => n415);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => n768,
                           QN => n416);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => n353
                           , QN => n417);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => n354
                           , QN => n418);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => n355
                           , QN => n419);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3195, CK => CLK, Q => n356
                           , QN => n420);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3194, CK => CLK, Q => n357
                           , QN => n421);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3193, CK => CLK, Q => n358
                           , QN => n422);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3192, CK => CLK, Q => n359
                           , QN => n423);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3191, CK => CLK, Q => n360
                           , QN => n424);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3190, CK => CLK, Q => n361
                           , QN => n425);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3189, CK => CLK, Q => n362
                           , QN => n426);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3188, CK => CLK, Q => n363
                           , QN => n427);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3187, CK => CLK, Q => n364
                           , QN => n428);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3186, CK => CLK, Q => n365
                           , QN => n429);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3185, CK => CLK, Q => n366
                           , QN => n430);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3184, CK => CLK, Q => n367
                           , QN => n431);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3183, CK => CLK, Q => n368
                           , QN => n432);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3182, CK => CLK, Q => n369
                           , QN => n433);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3181, CK => CLK, Q => n370
                           , QN => n434);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3180, CK => CLK, Q => n371
                           , QN => n435);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3179, CK => CLK, Q => n372
                           , QN => n436);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3178, CK => CLK, Q => n373
                           , QN => n437);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3177, CK => CLK, Q => n374
                           , QN => n438);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3176, CK => CLK, Q => n375,
                           QN => n439);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3175, CK => CLK, Q => n376,
                           QN => n440);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3174, CK => CLK, Q => n377,
                           QN => n441);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3173, CK => CLK, Q => n378,
                           QN => n442);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3172, CK => CLK, Q => n379,
                           QN => n443);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3171, CK => CLK, Q => n380,
                           QN => n444);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3170, CK => CLK, Q => n381,
                           QN => n445);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3169, CK => CLK, Q => n382,
                           QN => n446);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3168, CK => CLK, Q => n383,
                           QN => n447);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3167, CK => CLK, Q => n384,
                           QN => n448);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3166, CK => CLK, Q => 
                           n3956, QN => n_1236);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3165, CK => CLK, Q => 
                           n3955, QN => n_1237);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3164, CK => CLK, Q => 
                           n3954, QN => n_1238);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3163, CK => CLK, Q => 
                           n3953, QN => n_1239);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3162, CK => CLK, Q => 
                           n3952, QN => n_1240);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3161, CK => CLK, Q => 
                           n3951, QN => n_1241);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3160, CK => CLK, Q => 
                           n3950, QN => n_1242);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3159, CK => CLK, Q => 
                           n3949, QN => n_1243);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3158, CK => CLK, Q => 
                           n3948, QN => n_1244);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3157, CK => CLK, Q => 
                           n3947, QN => n_1245);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3156, CK => CLK, Q => 
                           n3946, QN => n_1246);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3155, CK => CLK, Q => 
                           n3945, QN => n_1247);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3154, CK => CLK, Q => 
                           n3944, QN => n_1248);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3153, CK => CLK, Q => 
                           n3943, QN => n_1249);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3152, CK => CLK, Q => 
                           n3942, QN => n_1250);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3151, CK => CLK, Q => 
                           n3941, QN => n_1251);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3150, CK => CLK, Q => 
                           n3940, QN => n_1252);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3149, CK => CLK, Q => 
                           n3939, QN => n_1253);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3148, CK => CLK, Q => 
                           n3938, QN => n_1254);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3147, CK => CLK, Q => 
                           n3937, QN => n_1255);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3146, CK => CLK, Q => 
                           n3936, QN => n_1256);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3145, CK => CLK, Q => 
                           n3935, QN => n_1257);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3144, CK => CLK, Q => n3934
                           , QN => n_1258);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3143, CK => CLK, Q => n3933
                           , QN => n_1259);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3142, CK => CLK, Q => n3932
                           , QN => n_1260);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3141, CK => CLK, Q => n3931
                           , QN => n_1261);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3140, CK => CLK, Q => n3930
                           , QN => n_1262);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3139, CK => CLK, Q => n3929
                           , QN => n_1263);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3138, CK => CLK, Q => n3928
                           , QN => n_1264);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3137, CK => CLK, Q => n3927
                           , QN => n_1265);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3136, CK => CLK, Q => n3926
                           , QN => n_1266);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3135, CK => CLK, Q => n3925
                           , QN => n_1267);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3134, CK => CLK, Q => 
                           n3924, QN => n_1268);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3133, CK => CLK, Q => 
                           n3923, QN => n_1269);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3132, CK => CLK, Q => 
                           n3922, QN => n_1270);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3131, CK => CLK, Q => 
                           n3921, QN => n_1271);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3130, CK => CLK, Q => 
                           n3920, QN => n_1272);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3129, CK => CLK, Q => 
                           n3919, QN => n_1273);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3128, CK => CLK, Q => 
                           n3918, QN => n_1274);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3127, CK => CLK, Q => 
                           n3917, QN => n_1275);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3126, CK => CLK, Q => 
                           n3916, QN => n_1276);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3125, CK => CLK, Q => 
                           n3915, QN => n_1277);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3124, CK => CLK, Q => 
                           n3914, QN => n_1278);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3123, CK => CLK, Q => 
                           n3913, QN => n_1279);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3122, CK => CLK, Q => 
                           n3912, QN => n_1280);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3121, CK => CLK, Q => 
                           n3911, QN => n_1281);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3120, CK => CLK, Q => 
                           n3910, QN => n_1282);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3119, CK => CLK, Q => 
                           n3909, QN => n_1283);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3118, CK => CLK, Q => 
                           n3908, QN => n_1284);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3117, CK => CLK, Q => 
                           n3907, QN => n_1285);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3116, CK => CLK, Q => 
                           n3906, QN => n_1286);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3115, CK => CLK, Q => 
                           n3905, QN => n_1287);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3114, CK => CLK, Q => 
                           n3904, QN => n_1288);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3113, CK => CLK, Q => 
                           n3903, QN => n_1289);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3112, CK => CLK, Q => n3902
                           , QN => n_1290);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3111, CK => CLK, Q => n3901
                           , QN => n_1291);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3110, CK => CLK, Q => n3900
                           , QN => n_1292);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3109, CK => CLK, Q => n3899
                           , QN => n_1293);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3108, CK => CLK, Q => n3898
                           , QN => n_1294);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3107, CK => CLK, Q => n3897
                           , QN => n_1295);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3106, CK => CLK, Q => n3896
                           , QN => n_1296);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3105, CK => CLK, Q => n3895
                           , QN => n_1297);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3104, CK => CLK, Q => n3894
                           , QN => n_1298);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3103, CK => CLK, Q => n3893
                           , QN => n_1299);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3102, CK => CLK, Q => n769
                           , QN => n513);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3101, CK => CLK, Q => n770
                           , QN => n514);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3100, CK => CLK, Q => n771
                           , QN => n515);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3099, CK => CLK, Q => n772
                           , QN => n516);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3098, CK => CLK, Q => n773
                           , QN => n517);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3097, CK => CLK, Q => n774
                           , QN => n518);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3096, CK => CLK, Q => n775
                           , QN => n519);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3095, CK => CLK, Q => n776
                           , QN => n520);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3094, CK => CLK, Q => n777
                           , QN => n521);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3093, CK => CLK, Q => n778
                           , QN => n522);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3092, CK => CLK, Q => n779
                           , QN => n523);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3091, CK => CLK, Q => n780
                           , QN => n524);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3090, CK => CLK, Q => n781
                           , QN => n525);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3089, CK => CLK, Q => n782
                           , QN => n526);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3088, CK => CLK, Q => n783
                           , QN => n527);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3087, CK => CLK, Q => n784
                           , QN => n528);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3086, CK => CLK, Q => n785
                           , QN => n529);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3085, CK => CLK, Q => n786
                           , QN => n530);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3084, CK => CLK, Q => n787
                           , QN => n531);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3083, CK => CLK, Q => n788
                           , QN => n532);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3082, CK => CLK, Q => n789
                           , QN => n533);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3081, CK => CLK, Q => n790
                           , QN => n534);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3080, CK => CLK, Q => n791,
                           QN => n535);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3079, CK => CLK, Q => n792,
                           QN => n536);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3078, CK => CLK, Q => n793,
                           QN => n537);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3077, CK => CLK, Q => n794,
                           QN => n538);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3076, CK => CLK, Q => n795,
                           QN => n539);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3075, CK => CLK, Q => n796,
                           QN => n540);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3074, CK => CLK, Q => n797,
                           QN => n541);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3073, CK => CLK, Q => n798,
                           QN => n542);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3072, CK => CLK, Q => n799,
                           QN => n543);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3071, CK => CLK, Q => n800,
                           QN => n544);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3070, CK => CLK, Q => n449
                           , QN => n545);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3069, CK => CLK, Q => n450
                           , QN => n546);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3068, CK => CLK, Q => n451
                           , QN => n547);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3067, CK => CLK, Q => n452
                           , QN => n548);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3066, CK => CLK, Q => n453
                           , QN => n549);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3065, CK => CLK, Q => n454
                           , QN => n550);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3064, CK => CLK, Q => n455
                           , QN => n551);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3063, CK => CLK, Q => n456
                           , QN => n552);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3062, CK => CLK, Q => n457
                           , QN => n553);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3061, CK => CLK, Q => n458
                           , QN => n554);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3060, CK => CLK, Q => n459
                           , QN => n555);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3059, CK => CLK, Q => n460
                           , QN => n556);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3058, CK => CLK, Q => n461
                           , QN => n557);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3057, CK => CLK, Q => n462
                           , QN => n558);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3056, CK => CLK, Q => n463
                           , QN => n559);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3055, CK => CLK, Q => n464
                           , QN => n560);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3054, CK => CLK, Q => n465
                           , QN => n561);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3053, CK => CLK, Q => n466
                           , QN => n562);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3052, CK => CLK, Q => n467
                           , QN => n563);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3051, CK => CLK, Q => n468
                           , QN => n564);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3050, CK => CLK, Q => n469
                           , QN => n565);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3049, CK => CLK, Q => n470
                           , QN => n566);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3048, CK => CLK, Q => n471,
                           QN => n567);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3047, CK => CLK, Q => n472,
                           QN => n568);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => n473,
                           QN => n569);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => n474,
                           QN => n570);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => n475,
                           QN => n571);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => n476,
                           QN => n572);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => n477,
                           QN => n573);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => n478,
                           QN => n574);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => n479,
                           QN => n575);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => n480,
                           QN => n576);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => 
                           n3892, QN => n_1300);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => 
                           n3891, QN => n_1301);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => 
                           n3890, QN => n_1302);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => 
                           n3889, QN => n_1303);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => 
                           n3888, QN => n_1304);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => 
                           n3887, QN => n_1305);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => 
                           n3886, QN => n_1306);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => 
                           n3885, QN => n_1307);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => 
                           n3884, QN => n_1308);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => 
                           n3883, QN => n_1309);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => 
                           n3882, QN => n_1310);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => 
                           n3881, QN => n_1311);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => 
                           n3880, QN => n_1312);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => 
                           n3879, QN => n_1313);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => 
                           n3878, QN => n_1314);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => 
                           n3877, QN => n_1315);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => 
                           n3876, QN => n_1316);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => 
                           n3875, QN => n_1317);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => 
                           n3874, QN => n_1318);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => 
                           n3873, QN => n_1319);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => 
                           n3872, QN => n_1320);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => 
                           n3871, QN => n_1321);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => n3870
                           , QN => n_1322);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => n3869
                           , QN => n_1323);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => n3868
                           , QN => n_1324);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => n3867
                           , QN => n_1325);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => n3866
                           , QN => n_1326);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => n3865
                           , QN => n_1327);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => n3864
                           , QN => n_1328);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => n3863
                           , QN => n_1329);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => n3862
                           , QN => n_1330);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => n3861
                           , QN => n_1331);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => 
                           n3860, QN => n_1332);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => 
                           n3859, QN => n_1333);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => 
                           n3858, QN => n_1334);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => 
                           n3857, QN => n_1335);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => 
                           n3856, QN => n_1336);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => 
                           n3855, QN => n_1337);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => 
                           n3854, QN => n_1338);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => 
                           n3853, QN => n_1339);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => 
                           n3852, QN => n_1340);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => 
                           n3851, QN => n_1341);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => 
                           n3850, QN => n_1342);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => 
                           n3849, QN => n_1343);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => 
                           n3848, QN => n_1344);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => 
                           n3847, QN => n_1345);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => 
                           n3846, QN => n_1346);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => 
                           n3845, QN => n_1347);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => 
                           n3844, QN => n_1348);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => 
                           n3843, QN => n_1349);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => 
                           n3842, QN => n_1350);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => 
                           n3841, QN => n_1351);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => 
                           n3840, QN => n_1352);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => 
                           n3839, QN => n_1353);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => n3838
                           , QN => n_1354);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => n3837
                           , QN => n_1355);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n2982, CK => CLK, Q => n3836
                           , QN => n_1356);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n2981, CK => CLK, Q => n3835
                           , QN => n_1357);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n2980, CK => CLK, Q => n3834
                           , QN => n_1358);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n2979, CK => CLK, Q => n3833
                           , QN => n_1359);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n2978, CK => CLK, Q => n3832
                           , QN => n_1360);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n2977, CK => CLK, Q => n3831
                           , QN => n_1361);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n2976, CK => CLK, Q => n3830
                           , QN => n_1362);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n2975, CK => CLK, Q => n3829
                           , QN => n_1363);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n2974, CK => CLK, Q => n801
                           , QN => n641);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n2973, CK => CLK, Q => n802
                           , QN => n642);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n2972, CK => CLK, Q => n803
                           , QN => n643);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n2971, CK => CLK, Q => n804
                           , QN => n644);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n2970, CK => CLK, Q => n805
                           , QN => n645);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n2969, CK => CLK, Q => n806
                           , QN => n646);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n2968, CK => CLK, Q => n807
                           , QN => n647);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n2967, CK => CLK, Q => n808
                           , QN => n648);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n2966, CK => CLK, Q => n809
                           , QN => n649);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n2965, CK => CLK, Q => n810
                           , QN => n650);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n2964, CK => CLK, Q => n811
                           , QN => n651);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n2963, CK => CLK, Q => n812
                           , QN => n652);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n2962, CK => CLK, Q => n813
                           , QN => n653);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n2961, CK => CLK, Q => n814
                           , QN => n654);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n2960, CK => CLK, Q => n815
                           , QN => n655);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n2959, CK => CLK, Q => n816
                           , QN => n656);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n2958, CK => CLK, Q => n817
                           , QN => n657);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n2957, CK => CLK, Q => n818
                           , QN => n658);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n2956, CK => CLK, Q => n819
                           , QN => n659);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n2955, CK => CLK, Q => n820
                           , QN => n660);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n2954, CK => CLK, Q => n821
                           , QN => n661);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n2953, CK => CLK, Q => n822
                           , QN => n662);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n2952, CK => CLK, Q => n823,
                           QN => n663);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n2951, CK => CLK, Q => n824,
                           QN => n664);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n2950, CK => CLK, Q => n825,
                           QN => n665);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n2949, CK => CLK, Q => n826,
                           QN => n666);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n2948, CK => CLK, Q => n827,
                           QN => n667);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n2947, CK => CLK, Q => n828,
                           QN => n668);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n2946, CK => CLK, Q => n829,
                           QN => n669);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n2945, CK => CLK, Q => n830,
                           QN => n670);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n2944, CK => CLK, Q => n831,
                           QN => n671);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n2943, CK => CLK, Q => n832,
                           QN => n672);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n2942, CK => CLK, Q => n481
                           , QN => n673);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n2941, CK => CLK, Q => n482
                           , QN => n674);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n2940, CK => CLK, Q => n483
                           , QN => n675);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n2939, CK => CLK, Q => n484
                           , QN => n676);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n2938, CK => CLK, Q => n485
                           , QN => n677);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n2937, CK => CLK, Q => n486
                           , QN => n678);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n2936, CK => CLK, Q => n487
                           , QN => n679);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n2935, CK => CLK, Q => n488
                           , QN => n680);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n2934, CK => CLK, Q => n489
                           , QN => n681);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n2933, CK => CLK, Q => n490
                           , QN => n682);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n2932, CK => CLK, Q => n491
                           , QN => n683);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n2931, CK => CLK, Q => n492
                           , QN => n684);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n2930, CK => CLK, Q => n493
                           , QN => n685);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n2929, CK => CLK, Q => n494
                           , QN => n686);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n2928, CK => CLK, Q => n495
                           , QN => n687);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n2927, CK => CLK, Q => n496
                           , QN => n688);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n2926, CK => CLK, Q => n497
                           , QN => n689);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n2925, CK => CLK, Q => n498
                           , QN => n690);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n2924, CK => CLK, Q => n499
                           , QN => n691);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n2923, CK => CLK, Q => n500
                           , QN => n692);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n2922, CK => CLK, Q => n501
                           , QN => n693);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n2921, CK => CLK, Q => n502
                           , QN => n694);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n2920, CK => CLK, Q => n503,
                           QN => n695);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n2919, CK => CLK, Q => n504,
                           QN => n696);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n2918, CK => CLK, Q => n505,
                           QN => n697);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n2917, CK => CLK, Q => n506,
                           QN => n698);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n2916, CK => CLK, Q => n507,
                           QN => n699);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n2915, CK => CLK, Q => n508,
                           QN => n700);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n2914, CK => CLK, Q => n509,
                           QN => n701);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n2913, CK => CLK, Q => n510,
                           QN => n702);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n2912, CK => CLK, Q => n511,
                           QN => n703);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n2911, CK => CLK, Q => n512,
                           QN => n704);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n2910, CK => CLK, Q => 
                           n3828, QN => n_1364);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n2909, CK => CLK, Q => 
                           n3827, QN => n_1365);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n2908, CK => CLK, Q => 
                           n3826, QN => n_1366);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n2907, CK => CLK, Q => 
                           n3825, QN => n_1367);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n2906, CK => CLK, Q => 
                           n3824, QN => n_1368);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n2905, CK => CLK, Q => 
                           n3823, QN => n_1369);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n2904, CK => CLK, Q => 
                           n3822, QN => n_1370);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n2903, CK => CLK, Q => 
                           n3821, QN => n_1371);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n2902, CK => CLK, Q => 
                           n3820, QN => n_1372);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n2901, CK => CLK, Q => 
                           n3819, QN => n_1373);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n2900, CK => CLK, Q => 
                           n3818, QN => n_1374);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n2899, CK => CLK, Q => 
                           n3817, QN => n_1375);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n2898, CK => CLK, Q => 
                           n3816, QN => n_1376);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n2897, CK => CLK, Q => 
                           n3815, QN => n_1377);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n2896, CK => CLK, Q => 
                           n3814, QN => n_1378);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n2895, CK => CLK, Q => 
                           n3813, QN => n_1379);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n2894, CK => CLK, Q => 
                           n3812, QN => n_1380);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n2893, CK => CLK, Q => 
                           n3811, QN => n_1381);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n2892, CK => CLK, Q => 
                           n3810, QN => n_1382);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n2891, CK => CLK, Q => 
                           n3809, QN => n_1383);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n2890, CK => CLK, Q => 
                           n3808, QN => n_1384);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n2889, CK => CLK, Q => 
                           n3807, QN => n_1385);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n2888, CK => CLK, Q => n3806
                           , QN => n_1386);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n2887, CK => CLK, Q => n3805
                           , QN => n_1387);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n2886, CK => CLK, Q => n3804
                           , QN => n_1388);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n2885, CK => CLK, Q => n3803
                           , QN => n_1389);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n2884, CK => CLK, Q => n3802
                           , QN => n_1390);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n2883, CK => CLK, Q => n3801
                           , QN => n_1391);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n2882, CK => CLK, Q => n3800
                           , QN => n_1392);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n2881, CK => CLK, Q => n3799
                           , QN => n_1393);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n2880, CK => CLK, Q => n3798
                           , QN => n_1394);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n2879, CK => CLK, Q => n3797
                           , QN => n_1395);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n2878, CK => CLK, Q => 
                           n3796, QN => n_1396);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n2877, CK => CLK, Q => 
                           n3795, QN => n_1397);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n2876, CK => CLK, Q => 
                           n3794, QN => n_1398);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n2875, CK => CLK, Q => 
                           n3793, QN => n_1399);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n2874, CK => CLK, Q => 
                           n3792, QN => n_1400);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n2873, CK => CLK, Q => 
                           n3791, QN => n_1401);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n2872, CK => CLK, Q => 
                           n3790, QN => n_1402);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n2871, CK => CLK, Q => 
                           n3789, QN => n_1403);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n2870, CK => CLK, Q => 
                           n3788, QN => n_1404);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n2869, CK => CLK, Q => 
                           n3787, QN => n_1405);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n2868, CK => CLK, Q => 
                           n3786, QN => n_1406);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n2867, CK => CLK, Q => 
                           n3785, QN => n_1407);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n2866, CK => CLK, Q => 
                           n3784, QN => n_1408);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => 
                           n3783, QN => n_1409);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => 
                           n3782, QN => n_1410);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => 
                           n3781, QN => n_1411);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => 
                           n3780, QN => n_1412);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => 
                           n3779, QN => n_1413);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n2860, CK => CLK, Q => 
                           n3778, QN => n_1414);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n2859, CK => CLK, Q => 
                           n3777, QN => n_1415);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n2858, CK => CLK, Q => 
                           n3776, QN => n_1416);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n2857, CK => CLK, Q => 
                           n3775, QN => n_1417);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n2856, CK => CLK, Q => n3774
                           , QN => n_1418);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n2855, CK => CLK, Q => n3773
                           , QN => n_1419);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n2854, CK => CLK, Q => n3772
                           , QN => n_1420);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n2853, CK => CLK, Q => n3771
                           , QN => n_1421);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n2852, CK => CLK, Q => n3770
                           , QN => n_1422);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n2851, CK => CLK, Q => n3769
                           , QN => n_1423);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n2850, CK => CLK, Q => n3768
                           , QN => n_1424);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n2849, CK => CLK, Q => n3767
                           , QN => n_1425);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n2848, CK => CLK, Q => n3766
                           , QN => n_1426);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n2847, CK => CLK, Q => n3765
                           , QN => n_1427);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n2846, CK => CLK, Q => 
                           n3764, QN => n_1428);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n2845, CK => CLK, Q => 
                           n3763, QN => n_1429);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n2844, CK => CLK, Q => 
                           n3762, QN => n_1430);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n2843, CK => CLK, Q => 
                           n3761, QN => n_1431);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n2842, CK => CLK, Q => 
                           n3760, QN => n_1432);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n2841, CK => CLK, Q => 
                           n3759, QN => n_1433);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n2840, CK => CLK, Q => 
                           n3758, QN => n_1434);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => 
                           n3757, QN => n_1435);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n2838, CK => CLK, Q => 
                           n3756, QN => n_1436);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n2837, CK => CLK, Q => 
                           n3755, QN => n_1437);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n2836, CK => CLK, Q => 
                           n3754, QN => n_1438);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n2835, CK => CLK, Q => 
                           n3753, QN => n_1439);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n2834, CK => CLK, Q => 
                           n3752, QN => n_1440);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n2833, CK => CLK, Q => 
                           n3751, QN => n_1441);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n2832, CK => CLK, Q => 
                           n3750, QN => n_1442);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n2831, CK => CLK, Q => 
                           n3749, QN => n_1443);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n2830, CK => CLK, Q => 
                           n3748, QN => n_1444);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n2829, CK => CLK, Q => 
                           n3747, QN => n_1445);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n2828, CK => CLK, Q => 
                           n3746, QN => n_1446);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n2827, CK => CLK, Q => 
                           n3745, QN => n_1447);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n2826, CK => CLK, Q => 
                           n3744, QN => n_1448);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n2825, CK => CLK, Q => 
                           n3743, QN => n_1449);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n2824, CK => CLK, Q => n3742
                           , QN => n_1450);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n2823, CK => CLK, Q => n3741
                           , QN => n_1451);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n2822, CK => CLK, Q => n3740
                           , QN => n_1452);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n2821, CK => CLK, Q => n3739
                           , QN => n_1453);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n2820, CK => CLK, Q => n3738
                           , QN => n_1454);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n2819, CK => CLK, Q => n3737
                           , QN => n_1455);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n2818, CK => CLK, Q => n3736
                           , QN => n_1456);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n2817, CK => CLK, Q => n3735
                           , QN => n_1457);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n2816, CK => CLK, Q => n3734
                           , QN => n_1458);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n2815, CK => CLK, Q => n3733
                           , QN => n_1459);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n2814, CK => CLK, Q => 
                           n3732, QN => n_1460);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n2813, CK => CLK, Q => 
                           n3731, QN => n_1461);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n2812, CK => CLK, Q => 
                           n3730, QN => n_1462);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n2811, CK => CLK, Q => 
                           n3729, QN => n_1463);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n2810, CK => CLK, Q => 
                           n3728, QN => n_1464);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n2809, CK => CLK, Q => 
                           n3727, QN => n_1465);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n2808, CK => CLK, Q => 
                           n3726, QN => n_1466);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n2807, CK => CLK, Q => 
                           n3725, QN => n_1467);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n2806, CK => CLK, Q => 
                           n3724, QN => n_1468);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n2805, CK => CLK, Q => 
                           n3723, QN => n_1469);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n2804, CK => CLK, Q => 
                           n3722, QN => n_1470);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n2803, CK => CLK, Q => 
                           n3721, QN => n_1471);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n2802, CK => CLK, Q => 
                           n3720, QN => n_1472);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n2801, CK => CLK, Q => 
                           n3719, QN => n_1473);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n2800, CK => CLK, Q => 
                           n3718, QN => n_1474);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n2799, CK => CLK, Q => 
                           n3717, QN => n_1475);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n2798, CK => CLK, Q => 
                           n3716, QN => n_1476);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n2797, CK => CLK, Q => 
                           n3715, QN => n_1477);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n2796, CK => CLK, Q => 
                           n3714, QN => n_1478);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n2795, CK => CLK, Q => 
                           n3713, QN => n_1479);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n2794, CK => CLK, Q => 
                           n3712, QN => n_1480);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n2793, CK => CLK, Q => 
                           n3711, QN => n_1481);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n2792, CK => CLK, Q => n3710
                           , QN => n_1482);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n2791, CK => CLK, Q => n3709
                           , QN => n_1483);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n2790, CK => CLK, Q => n3708
                           , QN => n_1484);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n2789, CK => CLK, Q => n3707
                           , QN => n_1485);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n2788, CK => CLK, Q => n3706
                           , QN => n_1486);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n2787, CK => CLK, Q => n3705
                           , QN => n_1487);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n2786, CK => CLK, Q => n3704
                           , QN => n_1488);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n2785, CK => CLK, Q => n3703
                           , QN => n_1489);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n2784, CK => CLK, Q => n3702
                           , QN => n_1490);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n2783, CK => CLK, Q => n3701
                           , QN => n_1491);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n2782, CK => CLK, Q => n897
                           , QN => n833);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n2781, CK => CLK, Q => n898
                           , QN => n834);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n2780, CK => CLK, Q => n899
                           , QN => n835);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n2779, CK => CLK, Q => n900
                           , QN => n836);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n2778, CK => CLK, Q => n901
                           , QN => n837);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n2777, CK => CLK, Q => n902
                           , QN => n838);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n2776, CK => CLK, Q => n903
                           , QN => n839);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n2775, CK => CLK, Q => n904
                           , QN => n840);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n2774, CK => CLK, Q => n905
                           , QN => n841);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n2773, CK => CLK, Q => n906
                           , QN => n842);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n2772, CK => CLK, Q => n907
                           , QN => n843);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n2771, CK => CLK, Q => n908
                           , QN => n844);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n2770, CK => CLK, Q => n909
                           , QN => n845);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n2769, CK => CLK, Q => n910
                           , QN => n846);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n2768, CK => CLK, Q => n911
                           , QN => n847);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n2767, CK => CLK, Q => n912
                           , QN => n848);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n2766, CK => CLK, Q => n913
                           , QN => n849);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n2765, CK => CLK, Q => n914
                           , QN => n850);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n2764, CK => CLK, Q => n915
                           , QN => n851);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n2763, CK => CLK, Q => n916
                           , QN => n852);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n2762, CK => CLK, Q => n917
                           , QN => n853);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n2761, CK => CLK, Q => n918
                           , QN => n854);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n2760, CK => CLK, Q => n919,
                           QN => n855);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n2759, CK => CLK, Q => n920,
                           QN => n856);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n2758, CK => CLK, Q => n921,
                           QN => n857);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n2757, CK => CLK, Q => n922,
                           QN => n858);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n2756, CK => CLK, Q => n923,
                           QN => n859);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n2755, CK => CLK, Q => n924,
                           QN => n860);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n2754, CK => CLK, Q => n925,
                           QN => n861);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n2753, CK => CLK, Q => n926,
                           QN => n862);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n2752, CK => CLK, Q => n927,
                           QN => n863);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n2751, CK => CLK, Q => n928,
                           QN => n864);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n2750, CK => CLK, Q => n577
                           , QN => n865);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n2749, CK => CLK, Q => n578
                           , QN => n866);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n2748, CK => CLK, Q => n579
                           , QN => n867);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n2747, CK => CLK, Q => n580
                           , QN => n868);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n2746, CK => CLK, Q => n581
                           , QN => n869);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n2745, CK => CLK, Q => n582
                           , QN => n870);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n2744, CK => CLK, Q => n583
                           , QN => n871);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n2743, CK => CLK, Q => n584
                           , QN => n872);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n2742, CK => CLK, Q => n585
                           , QN => n873);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n2741, CK => CLK, Q => n586
                           , QN => n874);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n2740, CK => CLK, Q => n587
                           , QN => n875);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n2739, CK => CLK, Q => n588
                           , QN => n876);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n2738, CK => CLK, Q => n589
                           , QN => n877);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n2737, CK => CLK, Q => n590
                           , QN => n878);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n2736, CK => CLK, Q => n591
                           , QN => n879);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n2735, CK => CLK, Q => n592
                           , QN => n880);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n2734, CK => CLK, Q => n593
                           , QN => n881);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n2733, CK => CLK, Q => n594
                           , QN => n882);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n2732, CK => CLK, Q => n595
                           , QN => n883);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n2731, CK => CLK, Q => n596
                           , QN => n884);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n2730, CK => CLK, Q => n597
                           , QN => n885);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n2729, CK => CLK, Q => n598
                           , QN => n886);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n2728, CK => CLK, Q => n599,
                           QN => n887);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n2727, CK => CLK, Q => n600,
                           QN => n888);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n2726, CK => CLK, Q => n601,
                           QN => n889);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n2725, CK => CLK, Q => n602,
                           QN => n890);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n2724, CK => CLK, Q => n603,
                           QN => n891);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n2723, CK => CLK, Q => n604,
                           QN => n892);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n2722, CK => CLK, Q => n605,
                           QN => n893);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n2721, CK => CLK, Q => n606,
                           QN => n894);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n2720, CK => CLK, Q => n607,
                           QN => n895);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n2719, CK => CLK, Q => n608,
                           QN => n896);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n2718, CK => CLK, Q => 
                           n3700, QN => n_1492);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n2717, CK => CLK, Q => 
                           n3699, QN => n_1493);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n2716, CK => CLK, Q => 
                           n3698, QN => n_1494);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n2715, CK => CLK, Q => 
                           n3697, QN => n_1495);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n2714, CK => CLK, Q => 
                           n3696, QN => n_1496);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n2713, CK => CLK, Q => 
                           n3695, QN => n_1497);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n2712, CK => CLK, Q => 
                           n3694, QN => n_1498);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n2711, CK => CLK, Q => 
                           n3693, QN => n_1499);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n2710, CK => CLK, Q => 
                           n3692, QN => n_1500);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n2709, CK => CLK, Q => 
                           n3691, QN => n_1501);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n2708, CK => CLK, Q => 
                           n3690, QN => n_1502);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n2707, CK => CLK, Q => 
                           n3689, QN => n_1503);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n2706, CK => CLK, Q => 
                           n3688, QN => n_1504);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n2705, CK => CLK, Q => 
                           n3687, QN => n_1505);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n2704, CK => CLK, Q => 
                           n3686, QN => n_1506);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n2703, CK => CLK, Q => 
                           n3685, QN => n_1507);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n2702, CK => CLK, Q => 
                           n3684, QN => n_1508);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n2701, CK => CLK, Q => 
                           n3683, QN => n_1509);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n2700, CK => CLK, Q => 
                           n3682, QN => n_1510);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n2699, CK => CLK, Q => 
                           n3681, QN => n_1511);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n2698, CK => CLK, Q => 
                           n3680, QN => n_1512);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n2697, CK => CLK, Q => 
                           n3679, QN => n_1513);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n2696, CK => CLK, Q => n3678
                           , QN => n_1514);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n2695, CK => CLK, Q => n3677
                           , QN => n_1515);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n2694, CK => CLK, Q => n3676
                           , QN => n_1516);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n2693, CK => CLK, Q => n3675
                           , QN => n_1517);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n2692, CK => CLK, Q => n3674
                           , QN => n_1518);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n2691, CK => CLK, Q => n3673
                           , QN => n_1519);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n2690, CK => CLK, Q => n3672
                           , QN => n_1520);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n2689, CK => CLK, Q => n3671
                           , QN => n_1521);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n2688, CK => CLK, Q => n3670
                           , QN => n_1522);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n2687, CK => CLK, Q => n3669
                           , QN => n_1523);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n2686, CK => CLK, Q => 
                           n3668, QN => n_1524);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n2685, CK => CLK, Q => 
                           n3667, QN => n_1525);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n2684, CK => CLK, Q => 
                           n3666, QN => n_1526);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n2683, CK => CLK, Q => 
                           n3665, QN => n_1527);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n2682, CK => CLK, Q => 
                           n3664, QN => n_1528);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n2681, CK => CLK, Q => 
                           n3663, QN => n_1529);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n2680, CK => CLK, Q => 
                           n3662, QN => n_1530);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n2679, CK => CLK, Q => 
                           n3661, QN => n_1531);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n2678, CK => CLK, Q => 
                           n3660, QN => n_1532);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n2677, CK => CLK, Q => 
                           n3659, QN => n_1533);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n2676, CK => CLK, Q => 
                           n3658, QN => n_1534);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n2675, CK => CLK, Q => 
                           n3657, QN => n_1535);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n2674, CK => CLK, Q => 
                           n3656, QN => n_1536);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n2673, CK => CLK, Q => 
                           n3655, QN => n_1537);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n2672, CK => CLK, Q => 
                           n3654, QN => n_1538);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n2671, CK => CLK, Q => 
                           n3653, QN => n_1539);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n2670, CK => CLK, Q => 
                           n3652, QN => n_1540);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n2669, CK => CLK, Q => 
                           n3651, QN => n_1541);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n2668, CK => CLK, Q => 
                           n3650, QN => n_1542);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n2667, CK => CLK, Q => 
                           n3649, QN => n_1543);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n2666, CK => CLK, Q => 
                           n3648, QN => n_1544);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n2665, CK => CLK, Q => 
                           n3647, QN => n_1545);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n2664, CK => CLK, Q => n3646
                           , QN => n_1546);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n2663, CK => CLK, Q => n3645
                           , QN => n_1547);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n2662, CK => CLK, Q => n3644
                           , QN => n_1548);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n2661, CK => CLK, Q => n3643
                           , QN => n_1549);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n2660, CK => CLK, Q => n3642
                           , QN => n_1550);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n2659, CK => CLK, Q => n3641
                           , QN => n_1551);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n2658, CK => CLK, Q => n3640
                           , QN => n_1552);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n2657, CK => CLK, Q => n3639
                           , QN => n_1553);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n2656, CK => CLK, Q => n3638
                           , QN => n_1554);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n2655, CK => CLK, Q => n3637
                           , QN => n_1555);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n2654, CK => CLK, Q => n929
                           , QN => n961);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n2653, CK => CLK, Q => n930
                           , QN => n962);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n2652, CK => CLK, Q => n931
                           , QN => n963);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n2651, CK => CLK, Q => n932
                           , QN => n964);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n2650, CK => CLK, Q => n933
                           , QN => n965);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n2649, CK => CLK, Q => n934
                           , QN => n966);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n2648, CK => CLK, Q => n935
                           , QN => n967);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n2647, CK => CLK, Q => n936
                           , QN => n968);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n2646, CK => CLK, Q => n937
                           , QN => n969);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n2645, CK => CLK, Q => n938
                           , QN => n970);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n2644, CK => CLK, Q => n939
                           , QN => n971);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n2643, CK => CLK, Q => n940
                           , QN => n972);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n2642, CK => CLK, Q => n941
                           , QN => n973);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n2641, CK => CLK, Q => n942
                           , QN => n974);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n2640, CK => CLK, Q => n943
                           , QN => n975);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n2639, CK => CLK, Q => n944
                           , QN => n976);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n2638, CK => CLK, Q => n945
                           , QN => n977);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n2637, CK => CLK, Q => n946
                           , QN => n978);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n2636, CK => CLK, Q => n947
                           , QN => n979);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n2635, CK => CLK, Q => n948
                           , QN => n980);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n2634, CK => CLK, Q => n949
                           , QN => n981);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n2633, CK => CLK, Q => n950
                           , QN => n982);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n2632, CK => CLK, Q => n951,
                           QN => n983);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n2631, CK => CLK, Q => n952,
                           QN => n984);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n2630, CK => CLK, Q => n953,
                           QN => n985);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n2629, CK => CLK, Q => n954,
                           QN => n986);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n2628, CK => CLK, Q => n955,
                           QN => n987);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n2627, CK => CLK, Q => n956,
                           QN => n988);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n2626, CK => CLK, Q => n957,
                           QN => n989);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n2625, CK => CLK, Q => n958,
                           QN => n990);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n2624, CK => CLK, Q => n959,
                           QN => n991);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n2623, CK => CLK, Q => n960,
                           QN => n992);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n2622, CK => CLK, Q => n609
                           , QN => n993);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n2621, CK => CLK, Q => n610
                           , QN => n994);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n2620, CK => CLK, Q => n611
                           , QN => n995);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n2619, CK => CLK, Q => n612
                           , QN => n996);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n2618, CK => CLK, Q => n613
                           , QN => n997);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n2617, CK => CLK, Q => n614
                           , QN => n998);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n2616, CK => CLK, Q => n615
                           , QN => n999);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n2615, CK => CLK, Q => n616
                           , QN => n1000);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n2614, CK => CLK, Q => n617
                           , QN => n1001);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n2613, CK => CLK, Q => n618
                           , QN => n1002);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n2612, CK => CLK, Q => n619
                           , QN => n1003);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n2611, CK => CLK, Q => n620
                           , QN => n1004);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n2610, CK => CLK, Q => n621
                           , QN => n1005);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n2609, CK => CLK, Q => n622
                           , QN => n1006);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n2608, CK => CLK, Q => n623
                           , QN => n1007);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n2607, CK => CLK, Q => n624
                           , QN => n1008);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n2606, CK => CLK, Q => n625
                           , QN => n1009);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n2605, CK => CLK, Q => n626
                           , QN => n1010);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n2604, CK => CLK, Q => n627
                           , QN => n1011);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n2603, CK => CLK, Q => n628
                           , QN => n1012);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n2602, CK => CLK, Q => n629
                           , QN => n1013);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n2601, CK => CLK, Q => n630
                           , QN => n1014);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n2600, CK => CLK, Q => n631,
                           QN => n1015);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n2599, CK => CLK, Q => n632,
                           QN => n1016);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n2598, CK => CLK, Q => n633,
                           QN => n1017);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n2597, CK => CLK, Q => n634,
                           QN => n1018);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n2596, CK => CLK, Q => n635,
                           QN => n1019);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n2595, CK => CLK, Q => n636,
                           QN => n1020);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n2594, CK => CLK, Q => n637,
                           QN => n1021);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n2593, CK => CLK, Q => n638,
                           QN => n1022);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n2592, CK => CLK, Q => n639,
                           QN => n1023);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n2591, CK => CLK, Q => n640,
                           QN => n1024);
   OUT1_reg_31_inst : DFF_X1 port map( D => n2590, CK => CLK, Q => OUT1(31), QN
                           => n3636);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2589, CK => CLK, Q => OUT1(30), QN
                           => n3635);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2588, CK => CLK, Q => OUT1(29), QN
                           => n3634);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2587, CK => CLK, Q => OUT1(28), QN
                           => n3633);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2586, CK => CLK, Q => OUT1(27), QN
                           => n3632);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2585, CK => CLK, Q => OUT1(26), QN
                           => n3631);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2584, CK => CLK, Q => OUT1(25), QN
                           => n3630);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2583, CK => CLK, Q => OUT1(24), QN
                           => n3629);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2582, CK => CLK, Q => OUT1(23), QN
                           => n3628);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2581, CK => CLK, Q => OUT1(22), QN
                           => n3627);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2580, CK => CLK, Q => OUT1(21), QN
                           => n3626);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2579, CK => CLK, Q => OUT1(20), QN
                           => n3625);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2578, CK => CLK, Q => OUT1(19), QN
                           => n3624);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2577, CK => CLK, Q => OUT1(18), QN
                           => n3623);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2576, CK => CLK, Q => OUT1(17), QN
                           => n3622);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2575, CK => CLK, Q => OUT1(16), QN
                           => n3621);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2574, CK => CLK, Q => OUT1(15), QN
                           => n3620);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2573, CK => CLK, Q => OUT1(14), QN
                           => n3619);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2572, CK => CLK, Q => OUT1(13), QN
                           => n3618);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2571, CK => CLK, Q => OUT1(12), QN
                           => n3617);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2570, CK => CLK, Q => OUT1(11), QN
                           => n3616);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => OUT1(10), QN
                           => n3615);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => OUT1(9), QN 
                           => n2526);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => OUT1(8), QN 
                           => n2525);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => OUT1(7), QN 
                           => n2524);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => OUT1(6), QN 
                           => n2523);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => OUT1(5), QN 
                           => n2522);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => OUT1(4), QN 
                           => n2521);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => OUT1(3), QN 
                           => n2520);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => OUT1(2), QN 
                           => n2519);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => OUT1(1), QN 
                           => n2518);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => OUT1(0), QN 
                           => n2517);
   OUT2_reg_31_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => OUT2(31), QN
                           => n2516);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => OUT2(30), QN
                           => n2515);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => OUT2(29), QN
                           => n2514);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => OUT2(28), QN
                           => n2513);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => OUT2(27), QN
                           => n2512);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => OUT2(26), QN
                           => n2511);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => OUT2(25), QN
                           => n2510);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => OUT2(24), QN
                           => n2509);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => OUT2(23), QN
                           => n2508);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => OUT2(22), QN
                           => n2507);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => OUT2(21), QN
                           => n2506);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => OUT2(20), QN
                           => n2505);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => OUT2(19), QN
                           => n2504);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => OUT2(18), QN
                           => n2503);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => OUT2(17), QN
                           => n2502);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => OUT2(16), QN
                           => n2501);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => OUT2(15), QN
                           => n2500);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => OUT2(14), QN
                           => n2499);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => OUT2(13), QN
                           => n2498);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => OUT2(12), QN
                           => n2497);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => OUT2(11), QN
                           => n2496);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => OUT2(10), QN
                           => n2495);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => OUT2(9), QN 
                           => n2494);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => OUT2(8), QN 
                           => n2493);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => OUT2(7), QN 
                           => n2492);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => OUT2(6), QN 
                           => n2491);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => OUT2(5), QN 
                           => n2490);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => OUT2(4), QN 
                           => n2489);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => OUT2(3), QN 
                           => n2488);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => OUT2(2), QN 
                           => n2487);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => OUT2(1), QN 
                           => n2486);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2527, CK => CLK, Q => OUT2(0), QN 
                           => n2485);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1170, ZN => n1172);
   U4 : NAND2_X2 port map( A1 => RST, A2 => n1828, ZN => n1830);
   U5 : INV_X1 port map( A => n1153, ZN => n1025);
   U6 : INV_X2 port map( A => n1025, ZN => n1026);
   U7 : INV_X1 port map( A => n1154, ZN => n1027);
   U8 : INV_X2 port map( A => n1027, ZN => n1028);
   U9 : INV_X1 port map( A => n1155, ZN => n1029);
   U10 : INV_X2 port map( A => n1029, ZN => n1030);
   U11 : INV_X1 port map( A => n1156, ZN => n1031);
   U12 : INV_X2 port map( A => n1031, ZN => n1032);
   U13 : INV_X1 port map( A => n1157, ZN => n1033);
   U14 : INV_X2 port map( A => n1033, ZN => n1034);
   U15 : INV_X1 port map( A => n1158, ZN => n1035);
   U16 : INV_X2 port map( A => n1035, ZN => n1036);
   U17 : INV_X1 port map( A => n1163, ZN => n1037);
   U18 : INV_X2 port map( A => n1037, ZN => n1038);
   U19 : INV_X1 port map( A => n1164, ZN => n1039);
   U20 : INV_X2 port map( A => n1039, ZN => n1040);
   U21 : INV_X1 port map( A => n1165, ZN => n1041);
   U22 : INV_X2 port map( A => n1041, ZN => n1042);
   U23 : INV_X1 port map( A => n1166, ZN => n1043);
   U24 : INV_X2 port map( A => n1043, ZN => n1044);
   U25 : INV_X1 port map( A => n1167, ZN => n1045);
   U26 : INV_X2 port map( A => n1045, ZN => n1046);
   U27 : INV_X1 port map( A => n1168, ZN => n1047);
   U28 : INV_X2 port map( A => n1047, ZN => n1048);
   U29 : INV_X1 port map( A => n1169, ZN => n1049);
   U30 : INV_X2 port map( A => n1049, ZN => n1050);
   U31 : INV_X1 port map( A => n1151, ZN => n1051);
   U32 : INV_X2 port map( A => n1051, ZN => n1052);
   U33 : INV_X1 port map( A => n1152, ZN => n1053);
   U34 : INV_X2 port map( A => n1053, ZN => n1054);
   U35 : INV_X1 port map( A => n1148, ZN => n1055);
   U36 : INV_X2 port map( A => n1055, ZN => n1056);
   U37 : INV_X1 port map( A => n1149, ZN => n1057);
   U38 : INV_X2 port map( A => n1057, ZN => n1058);
   U39 : INV_X1 port map( A => n1146, ZN => n1059);
   U40 : INV_X2 port map( A => n1059, ZN => n1060);
   U41 : INV_X1 port map( A => n1147, ZN => n1061);
   U42 : INV_X2 port map( A => n1061, ZN => n1062);
   U43 : INV_X1 port map( A => n1144, ZN => n1063);
   U44 : INV_X2 port map( A => n1063, ZN => n1064);
   U45 : INV_X1 port map( A => n1145, ZN => n1065);
   U46 : INV_X2 port map( A => n1065, ZN => n1066);
   U47 : INV_X1 port map( A => n1142, ZN => n1067);
   U48 : INV_X2 port map( A => n1067, ZN => n1068);
   U49 : INV_X1 port map( A => n1143, ZN => n1069);
   U50 : INV_X2 port map( A => n1069, ZN => n1070);
   U51 : INV_X1 port map( A => n1136, ZN => n1071);
   U52 : INV_X2 port map( A => n1071, ZN => n1072);
   U53 : INV_X1 port map( A => n1140, ZN => n1073);
   U54 : INV_X2 port map( A => n1073, ZN => n1074);
   U55 : INV_X1 port map( A => n1132, ZN => n1075);
   U56 : INV_X2 port map( A => n1075, ZN => n1076);
   U57 : INV_X1 port map( A => n1134, ZN => n1077);
   U58 : INV_X2 port map( A => n1077, ZN => n1078);
   U59 : INV_X1 port map( A => n1128, ZN => n1079);
   U60 : INV_X2 port map( A => n1079, ZN => n1080);
   U61 : INV_X1 port map( A => n1130, ZN => n1081);
   U62 : INV_X2 port map( A => n1081, ZN => n1082);
   U63 : INV_X1 port map( A => n1124, ZN => n1083);
   U64 : INV_X2 port map( A => n1083, ZN => n1084);
   U65 : INV_X1 port map( A => n1126, ZN => n1085);
   U66 : INV_X2 port map( A => n1085, ZN => n1086);
   U67 : INV_X1 port map( A => n1090, ZN => n1087);
   U68 : INV_X2 port map( A => n1087, ZN => n1088);
   U69 : AND2_X2 port map( A1 => n1811, A2 => n1802, ZN => n1189);
   U70 : AND2_X2 port map( A1 => n1803, A2 => n1804, ZN => n1179);
   U71 : AND2_X2 port map( A1 => n1806, A2 => n1820, ZN => n1208);
   U72 : AND2_X2 port map( A1 => n2469, A2 => n2460, ZN => n1847);
   U73 : AND2_X2 port map( A1 => n2461, A2 => n2462, ZN => n1837);
   U74 : AND2_X2 port map( A1 => n2464, A2 => n2478, ZN => n1866);
   U75 : AND2_X2 port map( A1 => n1824, A2 => n1807, ZN => n1218);
   U76 : AND2_X2 port map( A1 => n2482, A2 => n2465, ZN => n1876);
   U77 : AND2_X2 port map( A1 => n1811, A2 => n1806, ZN => n1194);
   U78 : AND2_X2 port map( A1 => n1803, A2 => n1807, ZN => n1184);
   U79 : AND2_X2 port map( A1 => n1802, A2 => n1820, ZN => n1203);
   U80 : AND2_X2 port map( A1 => n2469, A2 => n2464, ZN => n1852);
   U81 : AND2_X2 port map( A1 => n2461, A2 => n2465, ZN => n1842);
   U82 : AND2_X2 port map( A1 => n2460, A2 => n2478, ZN => n1861);
   U83 : AND2_X2 port map( A1 => n1824, A2 => n1804, ZN => n1213);
   U84 : AND2_X2 port map( A1 => n2482, A2 => n2462, ZN => n1871);
   U85 : NAND2_X2 port map( A1 => n1811, A2 => n1804, ZN => n1192);
   U86 : NAND2_X2 port map( A1 => n1803, A2 => n1802, ZN => n1182);
   U87 : NAND2_X2 port map( A1 => n1807, A2 => n1820, ZN => n1211);
   U88 : NAND2_X2 port map( A1 => n2469, A2 => n2462, ZN => n1850);
   U89 : NAND2_X2 port map( A1 => n2461, A2 => n2460, ZN => n1840);
   U90 : NAND2_X2 port map( A1 => n2465, A2 => n2478, ZN => n1869);
   U91 : NAND2_X2 port map( A1 => n1824, A2 => n1806, ZN => n1221);
   U92 : NAND2_X2 port map( A1 => n2482, A2 => n2464, ZN => n1879);
   U93 : NAND2_X2 port map( A1 => n1811, A2 => n1807, ZN => n1197);
   U94 : NAND2_X2 port map( A1 => n1803, A2 => n1806, ZN => n1187);
   U95 : NAND2_X2 port map( A1 => n1804, A2 => n1820, ZN => n1206);
   U96 : NAND2_X2 port map( A1 => n2469, A2 => n2465, ZN => n1855);
   U97 : NAND2_X2 port map( A1 => n2461, A2 => n2464, ZN => n1845);
   U98 : NAND2_X2 port map( A1 => n2462, A2 => n2478, ZN => n1864);
   U99 : NAND2_X2 port map( A1 => n1824, A2 => n1802, ZN => n1216);
   U100 : NAND2_X2 port map( A1 => n2482, A2 => n2460, ZN => n1874);
   U101 : AND2_X2 port map( A1 => n1810, A2 => n1802, ZN => n1190);
   U102 : AND2_X2 port map( A1 => n1801, A2 => n1804, ZN => n1180);
   U103 : AND2_X2 port map( A1 => n1806, A2 => n1819, ZN => n1209);
   U104 : AND2_X2 port map( A1 => n2468, A2 => n2460, ZN => n1848);
   U105 : AND2_X2 port map( A1 => n2459, A2 => n2462, ZN => n1838);
   U106 : AND2_X2 port map( A1 => n2464, A2 => n2477, ZN => n1867);
   U107 : AND2_X2 port map( A1 => n1823, A2 => n1807, ZN => n1219);
   U108 : AND2_X2 port map( A1 => n2481, A2 => n2465, ZN => n1877);
   U109 : AND2_X2 port map( A1 => n1810, A2 => n1806, ZN => n1195);
   U110 : AND2_X2 port map( A1 => n1801, A2 => n1807, ZN => n1185);
   U111 : AND2_X2 port map( A1 => n1819, A2 => n1802, ZN => n1204);
   U112 : AND2_X2 port map( A1 => n2468, A2 => n2464, ZN => n1853);
   U113 : AND2_X2 port map( A1 => n2459, A2 => n2465, ZN => n1843);
   U114 : AND2_X2 port map( A1 => n2477, A2 => n2460, ZN => n1862);
   U115 : AND2_X2 port map( A1 => n1823, A2 => n1804, ZN => n1214);
   U116 : AND2_X2 port map( A1 => n2481, A2 => n2462, ZN => n1872);
   U117 : NAND2_X2 port map( A1 => n1810, A2 => n1804, ZN => n1193);
   U118 : NAND2_X2 port map( A1 => n1801, A2 => n1802, ZN => n1183);
   U119 : NAND2_X2 port map( A1 => n1807, A2 => n1819, ZN => n1212);
   U120 : NAND2_X2 port map( A1 => n2468, A2 => n2462, ZN => n1851);
   U121 : NAND2_X2 port map( A1 => n2459, A2 => n2460, ZN => n1841);
   U122 : NAND2_X2 port map( A1 => n2465, A2 => n2477, ZN => n1870);
   U123 : NAND2_X2 port map( A1 => n1823, A2 => n1806, ZN => n1222);
   U124 : NAND2_X2 port map( A1 => n2481, A2 => n2464, ZN => n1880);
   U125 : OR2_X2 port map( A1 => RD1, A2 => n1827, ZN => n1170);
   U126 : NAND2_X2 port map( A1 => n1810, A2 => n1807, ZN => n1198);
   U127 : NAND2_X2 port map( A1 => n1801, A2 => n1806, ZN => n1188);
   U128 : NAND2_X2 port map( A1 => n1804, A2 => n1819, ZN => n1207);
   U129 : NAND2_X2 port map( A1 => n2468, A2 => n2465, ZN => n1856);
   U130 : NAND2_X2 port map( A1 => n2459, A2 => n2464, ZN => n1846);
   U131 : NAND2_X2 port map( A1 => n2462, A2 => n2477, ZN => n1865);
   U132 : NAND2_X2 port map( A1 => n1823, A2 => n1802, ZN => n1217);
   U133 : NAND2_X2 port map( A1 => n2481, A2 => n2460, ZN => n1875);
   U134 : OR2_X2 port map( A1 => RD2, A2 => n1827, ZN => n1828);
   U135 : MUX2_X1 port map( A => n130, B => n1089, S => n1088, Z => n3614);
   U136 : MUX2_X1 port map( A => n132, B => n1091, S => n1088, Z => n3613);
   U137 : MUX2_X1 port map( A => n134, B => n1092, S => n1088, Z => n3612);
   U138 : MUX2_X1 port map( A => n136, B => n1093, S => n1088, Z => n3611);
   U139 : MUX2_X1 port map( A => n138, B => n1094, S => n1088, Z => n3610);
   U140 : MUX2_X1 port map( A => n140, B => n1095, S => n1088, Z => n3609);
   U141 : MUX2_X1 port map( A => n142, B => n1096, S => n1088, Z => n3608);
   U142 : MUX2_X1 port map( A => n144, B => n1097, S => n1088, Z => n3607);
   U143 : MUX2_X1 port map( A => n146, B => n1098, S => n1088, Z => n3606);
   U144 : MUX2_X1 port map( A => n148, B => n1099, S => n1088, Z => n3605);
   U145 : MUX2_X1 port map( A => n150, B => n1100, S => n1088, Z => n3604);
   U146 : MUX2_X1 port map( A => n152, B => n1101, S => n1088, Z => n3603);
   U147 : MUX2_X1 port map( A => n154, B => n1102, S => n1088, Z => n3602);
   U148 : MUX2_X1 port map( A => n156, B => n1103, S => n1088, Z => n3601);
   U149 : MUX2_X1 port map( A => n158, B => n1104, S => n1088, Z => n3600);
   U150 : MUX2_X1 port map( A => n160, B => n1105, S => n1088, Z => n3599);
   U151 : MUX2_X1 port map( A => n162, B => n1106, S => n1088, Z => n3598);
   U152 : MUX2_X1 port map( A => n164, B => n1107, S => n1088, Z => n3597);
   U153 : MUX2_X1 port map( A => n166, B => n1108, S => n1088, Z => n3596);
   U154 : MUX2_X1 port map( A => n168, B => n1109, S => n1088, Z => n3595);
   U155 : MUX2_X1 port map( A => n170, B => n1110, S => n1088, Z => n3594);
   U156 : MUX2_X1 port map( A => n172, B => n1111, S => n1088, Z => n3593);
   U157 : MUX2_X1 port map( A => n174, B => n1112, S => n1088, Z => n3592);
   U158 : MUX2_X1 port map( A => n176, B => n1113, S => n1088, Z => n3591);
   U159 : MUX2_X1 port map( A => n178, B => n1114, S => n1088, Z => n3590);
   U160 : MUX2_X1 port map( A => n180, B => n1115, S => n1088, Z => n3589);
   U161 : MUX2_X1 port map( A => n182, B => n1116, S => n1088, Z => n3588);
   U162 : MUX2_X1 port map( A => n184, B => n1117, S => n1088, Z => n3587);
   U163 : MUX2_X1 port map( A => n186, B => n1118, S => n1088, Z => n3586);
   U164 : MUX2_X1 port map( A => n188, B => n1119, S => n1088, Z => n3585);
   U165 : MUX2_X1 port map( A => n190, B => n1120, S => n1088, Z => n3584);
   U166 : MUX2_X1 port map( A => n192, B => n1121, S => n1088, Z => n3583);
   U167 : OAI21_X1 port map( B1 => n1122, B2 => n1123, A => RST, ZN => n1090);
   U168 : MUX2_X1 port map( A => n2, B => n1089, S => n1084, Z => n3582);
   U169 : MUX2_X1 port map( A => n4, B => n1091, S => n1084, Z => n3581);
   U170 : MUX2_X1 port map( A => n6, B => n1092, S => n1084, Z => n3580);
   U171 : MUX2_X1 port map( A => n8, B => n1093, S => n1084, Z => n3579);
   U172 : MUX2_X1 port map( A => n10, B => n1094, S => n1084, Z => n3578);
   U173 : MUX2_X1 port map( A => n12, B => n1095, S => n1084, Z => n3577);
   U174 : MUX2_X1 port map( A => n14, B => n1096, S => n1084, Z => n3576);
   U175 : MUX2_X1 port map( A => n16, B => n1097, S => n1084, Z => n3575);
   U176 : MUX2_X1 port map( A => n18, B => n1098, S => n1084, Z => n3574);
   U177 : MUX2_X1 port map( A => n20, B => n1099, S => n1084, Z => n3573);
   U178 : MUX2_X1 port map( A => n22, B => n1100, S => n1084, Z => n3572);
   U179 : MUX2_X1 port map( A => n24, B => n1101, S => n1084, Z => n3571);
   U180 : MUX2_X1 port map( A => n26, B => n1102, S => n1084, Z => n3570);
   U181 : MUX2_X1 port map( A => n28, B => n1103, S => n1084, Z => n3569);
   U182 : MUX2_X1 port map( A => n30, B => n1104, S => n1084, Z => n3568);
   U183 : MUX2_X1 port map( A => n32, B => n1105, S => n1084, Z => n3567);
   U184 : MUX2_X1 port map( A => n34, B => n1106, S => n1084, Z => n3566);
   U185 : MUX2_X1 port map( A => n36, B => n1107, S => n1084, Z => n3565);
   U186 : MUX2_X1 port map( A => n38, B => n1108, S => n1084, Z => n3564);
   U187 : MUX2_X1 port map( A => n40, B => n1109, S => n1084, Z => n3563);
   U188 : MUX2_X1 port map( A => n42, B => n1110, S => n1084, Z => n3562);
   U189 : MUX2_X1 port map( A => n44, B => n1111, S => n1084, Z => n3561);
   U190 : MUX2_X1 port map( A => n46, B => n1112, S => n1084, Z => n3560);
   U191 : MUX2_X1 port map( A => n48, B => n1113, S => n1084, Z => n3559);
   U192 : MUX2_X1 port map( A => n50, B => n1114, S => n1084, Z => n3558);
   U193 : MUX2_X1 port map( A => n52, B => n1115, S => n1084, Z => n3557);
   U194 : MUX2_X1 port map( A => n54, B => n1116, S => n1084, Z => n3556);
   U195 : MUX2_X1 port map( A => n56, B => n1117, S => n1084, Z => n3555);
   U196 : MUX2_X1 port map( A => n58, B => n1118, S => n1084, Z => n3554);
   U197 : MUX2_X1 port map( A => n60, B => n1119, S => n1084, Z => n3553);
   U198 : MUX2_X1 port map( A => n62, B => n1120, S => n1084, Z => n3552);
   U199 : MUX2_X1 port map( A => n64, B => n1121, S => n1084, Z => n3551);
   U200 : OAI21_X1 port map( B1 => n1122, B2 => n1125, A => RST, ZN => n1124);
   U201 : MUX2_X1 port map( A => n4148, B => n1089, S => n1086, Z => n3550);
   U202 : MUX2_X1 port map( A => n4147, B => n1091, S => n1086, Z => n3549);
   U203 : MUX2_X1 port map( A => n4146, B => n1092, S => n1086, Z => n3548);
   U204 : MUX2_X1 port map( A => n4145, B => n1093, S => n1086, Z => n3547);
   U205 : MUX2_X1 port map( A => n4144, B => n1094, S => n1086, Z => n3546);
   U206 : MUX2_X1 port map( A => n4143, B => n1095, S => n1086, Z => n3545);
   U207 : MUX2_X1 port map( A => n4142, B => n1096, S => n1086, Z => n3544);
   U208 : MUX2_X1 port map( A => n4141, B => n1097, S => n1086, Z => n3543);
   U209 : MUX2_X1 port map( A => n4140, B => n1098, S => n1086, Z => n3542);
   U210 : MUX2_X1 port map( A => n4139, B => n1099, S => n1086, Z => n3541);
   U211 : MUX2_X1 port map( A => n4138, B => n1100, S => n1086, Z => n3540);
   U212 : MUX2_X1 port map( A => n4137, B => n1101, S => n1086, Z => n3539);
   U213 : MUX2_X1 port map( A => n4136, B => n1102, S => n1086, Z => n3538);
   U214 : MUX2_X1 port map( A => n4135, B => n1103, S => n1086, Z => n3537);
   U215 : MUX2_X1 port map( A => n4134, B => n1104, S => n1086, Z => n3536);
   U216 : MUX2_X1 port map( A => n4133, B => n1105, S => n1086, Z => n3535);
   U217 : MUX2_X1 port map( A => n4132, B => n1106, S => n1086, Z => n3534);
   U218 : MUX2_X1 port map( A => n4131, B => n1107, S => n1086, Z => n3533);
   U219 : MUX2_X1 port map( A => n4130, B => n1108, S => n1086, Z => n3532);
   U220 : MUX2_X1 port map( A => n4129, B => n1109, S => n1086, Z => n3531);
   U221 : MUX2_X1 port map( A => n4128, B => n1110, S => n1086, Z => n3530);
   U222 : MUX2_X1 port map( A => n4127, B => n1111, S => n1086, Z => n3529);
   U223 : MUX2_X1 port map( A => n4126, B => n1112, S => n1086, Z => n3528);
   U224 : MUX2_X1 port map( A => n4125, B => n1113, S => n1086, Z => n3527);
   U225 : MUX2_X1 port map( A => n4124, B => n1114, S => n1086, Z => n3526);
   U226 : MUX2_X1 port map( A => n4123, B => n1115, S => n1086, Z => n3525);
   U227 : MUX2_X1 port map( A => n4122, B => n1116, S => n1086, Z => n3524);
   U228 : MUX2_X1 port map( A => n4121, B => n1117, S => n1086, Z => n3523);
   U229 : MUX2_X1 port map( A => n4120, B => n1118, S => n1086, Z => n3522);
   U230 : MUX2_X1 port map( A => n4119, B => n1119, S => n1086, Z => n3521);
   U231 : MUX2_X1 port map( A => n4118, B => n1120, S => n1086, Z => n3520);
   U232 : MUX2_X1 port map( A => n4117, B => n1121, S => n1086, Z => n3519);
   U233 : OAI21_X1 port map( B1 => n1122, B2 => n1127, A => RST, ZN => n1126);
   U234 : MUX2_X1 port map( A => n4116, B => n1089, S => n1080, Z => n3518);
   U235 : MUX2_X1 port map( A => n4115, B => n1091, S => n1080, Z => n3517);
   U236 : MUX2_X1 port map( A => n4114, B => n1092, S => n1080, Z => n3516);
   U237 : MUX2_X1 port map( A => n4113, B => n1093, S => n1080, Z => n3515);
   U238 : MUX2_X1 port map( A => n4112, B => n1094, S => n1080, Z => n3514);
   U239 : MUX2_X1 port map( A => n4111, B => n1095, S => n1080, Z => n3513);
   U240 : MUX2_X1 port map( A => n4110, B => n1096, S => n1080, Z => n3512);
   U241 : MUX2_X1 port map( A => n4109, B => n1097, S => n1080, Z => n3511);
   U242 : MUX2_X1 port map( A => n4108, B => n1098, S => n1080, Z => n3510);
   U243 : MUX2_X1 port map( A => n4107, B => n1099, S => n1080, Z => n3509);
   U244 : MUX2_X1 port map( A => n4106, B => n1100, S => n1080, Z => n3508);
   U245 : MUX2_X1 port map( A => n4105, B => n1101, S => n1080, Z => n3507);
   U246 : MUX2_X1 port map( A => n4104, B => n1102, S => n1080, Z => n3506);
   U247 : MUX2_X1 port map( A => n4103, B => n1103, S => n1080, Z => n3505);
   U248 : MUX2_X1 port map( A => n4102, B => n1104, S => n1080, Z => n3504);
   U249 : MUX2_X1 port map( A => n4101, B => n1105, S => n1080, Z => n3503);
   U250 : MUX2_X1 port map( A => n4100, B => n1106, S => n1080, Z => n3502);
   U251 : MUX2_X1 port map( A => n4099, B => n1107, S => n1080, Z => n3501);
   U252 : MUX2_X1 port map( A => n4098, B => n1108, S => n1080, Z => n3500);
   U253 : MUX2_X1 port map( A => n4097, B => n1109, S => n1080, Z => n3499);
   U254 : MUX2_X1 port map( A => n4096, B => n1110, S => n1080, Z => n3498);
   U255 : MUX2_X1 port map( A => n4095, B => n1111, S => n1080, Z => n3497);
   U256 : MUX2_X1 port map( A => n4094, B => n1112, S => n1080, Z => n3496);
   U257 : MUX2_X1 port map( A => n4093, B => n1113, S => n1080, Z => n3495);
   U258 : MUX2_X1 port map( A => n4092, B => n1114, S => n1080, Z => n3494);
   U259 : MUX2_X1 port map( A => n4091, B => n1115, S => n1080, Z => n3493);
   U260 : MUX2_X1 port map( A => n4090, B => n1116, S => n1080, Z => n3492);
   U261 : MUX2_X1 port map( A => n4089, B => n1117, S => n1080, Z => n3491);
   U262 : MUX2_X1 port map( A => n4088, B => n1118, S => n1080, Z => n3490);
   U263 : MUX2_X1 port map( A => n4087, B => n1119, S => n1080, Z => n3489);
   U264 : MUX2_X1 port map( A => n4086, B => n1120, S => n1080, Z => n3488);
   U265 : MUX2_X1 port map( A => n4085, B => n1121, S => n1080, Z => n3487);
   U266 : OAI21_X1 port map( B1 => n1122, B2 => n1129, A => RST, ZN => n1128);
   U267 : MUX2_X1 port map( A => n129, B => n1089, S => n1082, Z => n3486);
   U268 : MUX2_X1 port map( A => n131, B => n1091, S => n1082, Z => n3485);
   U269 : MUX2_X1 port map( A => n133, B => n1092, S => n1082, Z => n3484);
   U270 : MUX2_X1 port map( A => n135, B => n1093, S => n1082, Z => n3483);
   U271 : MUX2_X1 port map( A => n137, B => n1094, S => n1082, Z => n3482);
   U272 : MUX2_X1 port map( A => n139, B => n1095, S => n1082, Z => n3481);
   U273 : MUX2_X1 port map( A => n141, B => n1096, S => n1082, Z => n3480);
   U274 : MUX2_X1 port map( A => n143, B => n1097, S => n1082, Z => n3479);
   U275 : MUX2_X1 port map( A => n145, B => n1098, S => n1082, Z => n3478);
   U276 : MUX2_X1 port map( A => n147, B => n1099, S => n1082, Z => n3477);
   U277 : MUX2_X1 port map( A => n149, B => n1100, S => n1082, Z => n3476);
   U278 : MUX2_X1 port map( A => n151, B => n1101, S => n1082, Z => n3475);
   U279 : MUX2_X1 port map( A => n153, B => n1102, S => n1082, Z => n3474);
   U280 : MUX2_X1 port map( A => n155, B => n1103, S => n1082, Z => n3473);
   U281 : MUX2_X1 port map( A => n157, B => n1104, S => n1082, Z => n3472);
   U282 : MUX2_X1 port map( A => n159, B => n1105, S => n1082, Z => n3471);
   U283 : MUX2_X1 port map( A => n161, B => n1106, S => n1082, Z => n3470);
   U284 : MUX2_X1 port map( A => n163, B => n1107, S => n1082, Z => n3469);
   U285 : MUX2_X1 port map( A => n165, B => n1108, S => n1082, Z => n3468);
   U286 : MUX2_X1 port map( A => n167, B => n1109, S => n1082, Z => n3467);
   U287 : MUX2_X1 port map( A => n169, B => n1110, S => n1082, Z => n3466);
   U288 : MUX2_X1 port map( A => n171, B => n1111, S => n1082, Z => n3465);
   U289 : MUX2_X1 port map( A => n173, B => n1112, S => n1082, Z => n3464);
   U290 : MUX2_X1 port map( A => n175, B => n1113, S => n1082, Z => n3463);
   U291 : MUX2_X1 port map( A => n177, B => n1114, S => n1082, Z => n3462);
   U292 : MUX2_X1 port map( A => n179, B => n1115, S => n1082, Z => n3461);
   U293 : MUX2_X1 port map( A => n181, B => n1116, S => n1082, Z => n3460);
   U294 : MUX2_X1 port map( A => n183, B => n1117, S => n1082, Z => n3459);
   U295 : MUX2_X1 port map( A => n185, B => n1118, S => n1082, Z => n3458);
   U296 : MUX2_X1 port map( A => n187, B => n1119, S => n1082, Z => n3457);
   U297 : MUX2_X1 port map( A => n189, B => n1120, S => n1082, Z => n3456);
   U298 : MUX2_X1 port map( A => n191, B => n1121, S => n1082, Z => n3455);
   U299 : OAI21_X1 port map( B1 => n1122, B2 => n1131, A => RST, ZN => n1130);
   U300 : MUX2_X1 port map( A => n1, B => n1089, S => n1076, Z => n3454);
   U301 : MUX2_X1 port map( A => n3, B => n1091, S => n1076, Z => n3453);
   U302 : MUX2_X1 port map( A => n5, B => n1092, S => n1076, Z => n3452);
   U303 : MUX2_X1 port map( A => n7, B => n1093, S => n1076, Z => n3451);
   U304 : MUX2_X1 port map( A => n9, B => n1094, S => n1076, Z => n3450);
   U305 : MUX2_X1 port map( A => n11, B => n1095, S => n1076, Z => n3449);
   U306 : MUX2_X1 port map( A => n13, B => n1096, S => n1076, Z => n3448);
   U307 : MUX2_X1 port map( A => n15, B => n1097, S => n1076, Z => n3447);
   U308 : MUX2_X1 port map( A => n17, B => n1098, S => n1076, Z => n3446);
   U309 : MUX2_X1 port map( A => n19, B => n1099, S => n1076, Z => n3445);
   U310 : MUX2_X1 port map( A => n21, B => n1100, S => n1076, Z => n3444);
   U311 : MUX2_X1 port map( A => n23, B => n1101, S => n1076, Z => n3443);
   U312 : MUX2_X1 port map( A => n25, B => n1102, S => n1076, Z => n3442);
   U313 : MUX2_X1 port map( A => n27, B => n1103, S => n1076, Z => n3441);
   U314 : MUX2_X1 port map( A => n29, B => n1104, S => n1076, Z => n3440);
   U315 : MUX2_X1 port map( A => n31, B => n1105, S => n1076, Z => n3439);
   U316 : MUX2_X1 port map( A => n33, B => n1106, S => n1076, Z => n3438);
   U317 : MUX2_X1 port map( A => n35, B => n1107, S => n1076, Z => n3437);
   U318 : MUX2_X1 port map( A => n37, B => n1108, S => n1076, Z => n3436);
   U319 : MUX2_X1 port map( A => n39, B => n1109, S => n1076, Z => n3435);
   U320 : MUX2_X1 port map( A => n41, B => n1110, S => n1076, Z => n3434);
   U321 : MUX2_X1 port map( A => n43, B => n1111, S => n1076, Z => n3433);
   U322 : MUX2_X1 port map( A => n45, B => n1112, S => n1076, Z => n3432);
   U323 : MUX2_X1 port map( A => n47, B => n1113, S => n1076, Z => n3431);
   U324 : MUX2_X1 port map( A => n49, B => n1114, S => n1076, Z => n3430);
   U325 : MUX2_X1 port map( A => n51, B => n1115, S => n1076, Z => n3429);
   U326 : MUX2_X1 port map( A => n53, B => n1116, S => n1076, Z => n3428);
   U327 : MUX2_X1 port map( A => n55, B => n1117, S => n1076, Z => n3427);
   U328 : MUX2_X1 port map( A => n57, B => n1118, S => n1076, Z => n3426);
   U329 : MUX2_X1 port map( A => n59, B => n1119, S => n1076, Z => n3425);
   U330 : MUX2_X1 port map( A => n61, B => n1120, S => n1076, Z => n3424);
   U331 : MUX2_X1 port map( A => n63, B => n1121, S => n1076, Z => n3423);
   U332 : OAI21_X1 port map( B1 => n1122, B2 => n1133, A => RST, ZN => n1132);
   U333 : MUX2_X1 port map( A => n4084, B => n1089, S => n1078, Z => n3422);
   U334 : MUX2_X1 port map( A => n4083, B => n1091, S => n1078, Z => n3421);
   U335 : MUX2_X1 port map( A => n4082, B => n1092, S => n1078, Z => n3420);
   U336 : MUX2_X1 port map( A => n4081, B => n1093, S => n1078, Z => n3419);
   U337 : MUX2_X1 port map( A => n4080, B => n1094, S => n1078, Z => n3418);
   U338 : MUX2_X1 port map( A => n4079, B => n1095, S => n1078, Z => n3417);
   U339 : MUX2_X1 port map( A => n4078, B => n1096, S => n1078, Z => n3416);
   U340 : MUX2_X1 port map( A => n4077, B => n1097, S => n1078, Z => n3415);
   U341 : MUX2_X1 port map( A => n4076, B => n1098, S => n1078, Z => n3414);
   U342 : MUX2_X1 port map( A => n4075, B => n1099, S => n1078, Z => n3413);
   U343 : MUX2_X1 port map( A => n4074, B => n1100, S => n1078, Z => n3412);
   U344 : MUX2_X1 port map( A => n4073, B => n1101, S => n1078, Z => n3411);
   U345 : MUX2_X1 port map( A => n4072, B => n1102, S => n1078, Z => n3410);
   U346 : MUX2_X1 port map( A => n4071, B => n1103, S => n1078, Z => n3409);
   U347 : MUX2_X1 port map( A => n4070, B => n1104, S => n1078, Z => n3408);
   U348 : MUX2_X1 port map( A => n4069, B => n1105, S => n1078, Z => n3407);
   U349 : MUX2_X1 port map( A => n4068, B => n1106, S => n1078, Z => n3406);
   U350 : MUX2_X1 port map( A => n4067, B => n1107, S => n1078, Z => n3405);
   U351 : MUX2_X1 port map( A => n4066, B => n1108, S => n1078, Z => n3404);
   U352 : MUX2_X1 port map( A => n4065, B => n1109, S => n1078, Z => n3403);
   U353 : MUX2_X1 port map( A => n4064, B => n1110, S => n1078, Z => n3402);
   U354 : MUX2_X1 port map( A => n4063, B => n1111, S => n1078, Z => n3401);
   U355 : MUX2_X1 port map( A => n4062, B => n1112, S => n1078, Z => n3400);
   U356 : MUX2_X1 port map( A => n4061, B => n1113, S => n1078, Z => n3399);
   U357 : MUX2_X1 port map( A => n4060, B => n1114, S => n1078, Z => n3398);
   U358 : MUX2_X1 port map( A => n4059, B => n1115, S => n1078, Z => n3397);
   U359 : MUX2_X1 port map( A => n4058, B => n1116, S => n1078, Z => n3396);
   U360 : MUX2_X1 port map( A => n4057, B => n1117, S => n1078, Z => n3395);
   U361 : MUX2_X1 port map( A => n4056, B => n1118, S => n1078, Z => n3394);
   U362 : MUX2_X1 port map( A => n4055, B => n1119, S => n1078, Z => n3393);
   U363 : MUX2_X1 port map( A => n4054, B => n1120, S => n1078, Z => n3392);
   U364 : MUX2_X1 port map( A => n4053, B => n1121, S => n1078, Z => n3391);
   U365 : OAI21_X1 port map( B1 => n1122, B2 => n1135, A => RST, ZN => n1134);
   U366 : MUX2_X1 port map( A => n4052, B => n1089, S => n1072, Z => n3390);
   U367 : MUX2_X1 port map( A => n4051, B => n1091, S => n1072, Z => n3389);
   U368 : MUX2_X1 port map( A => n4050, B => n1092, S => n1072, Z => n3388);
   U369 : MUX2_X1 port map( A => n4049, B => n1093, S => n1072, Z => n3387);
   U370 : MUX2_X1 port map( A => n4048, B => n1094, S => n1072, Z => n3386);
   U371 : MUX2_X1 port map( A => n4047, B => n1095, S => n1072, Z => n3385);
   U372 : MUX2_X1 port map( A => n4046, B => n1096, S => n1072, Z => n3384);
   U373 : MUX2_X1 port map( A => n4045, B => n1097, S => n1072, Z => n3383);
   U374 : MUX2_X1 port map( A => n4044, B => n1098, S => n1072, Z => n3382);
   U375 : MUX2_X1 port map( A => n4043, B => n1099, S => n1072, Z => n3381);
   U376 : MUX2_X1 port map( A => n4042, B => n1100, S => n1072, Z => n3380);
   U377 : MUX2_X1 port map( A => n4041, B => n1101, S => n1072, Z => n3379);
   U378 : MUX2_X1 port map( A => n4040, B => n1102, S => n1072, Z => n3378);
   U379 : MUX2_X1 port map( A => n4039, B => n1103, S => n1072, Z => n3377);
   U380 : MUX2_X1 port map( A => n4038, B => n1104, S => n1072, Z => n3376);
   U381 : MUX2_X1 port map( A => n4037, B => n1105, S => n1072, Z => n3375);
   U382 : MUX2_X1 port map( A => n4036, B => n1106, S => n1072, Z => n3374);
   U383 : MUX2_X1 port map( A => n4035, B => n1107, S => n1072, Z => n3373);
   U384 : MUX2_X1 port map( A => n4034, B => n1108, S => n1072, Z => n3372);
   U385 : MUX2_X1 port map( A => n4033, B => n1109, S => n1072, Z => n3371);
   U386 : MUX2_X1 port map( A => n4032, B => n1110, S => n1072, Z => n3370);
   U387 : MUX2_X1 port map( A => n4031, B => n1111, S => n1072, Z => n3369);
   U388 : MUX2_X1 port map( A => n4030, B => n1112, S => n1072, Z => n3368);
   U389 : MUX2_X1 port map( A => n4029, B => n1113, S => n1072, Z => n3367);
   U390 : MUX2_X1 port map( A => n4028, B => n1114, S => n1072, Z => n3366);
   U391 : MUX2_X1 port map( A => n4027, B => n1115, S => n1072, Z => n3365);
   U392 : MUX2_X1 port map( A => n4026, B => n1116, S => n1072, Z => n3364);
   U393 : MUX2_X1 port map( A => n4025, B => n1117, S => n1072, Z => n3363);
   U394 : MUX2_X1 port map( A => n4024, B => n1118, S => n1072, Z => n3362);
   U395 : MUX2_X1 port map( A => n4023, B => n1119, S => n1072, Z => n3361);
   U396 : MUX2_X1 port map( A => n4022, B => n1120, S => n1072, Z => n3360);
   U397 : MUX2_X1 port map( A => n4021, B => n1121, S => n1072, Z => n3359);
   U398 : OAI21_X1 port map( B1 => n1122, B2 => n1137, A => RST, ZN => n1136);
   U399 : NAND3_X1 port map( A1 => n1138, A2 => n1139, A3 => WR, ZN => n1122);
   U400 : MUX2_X1 port map( A => n705, B => n1089, S => n1074, Z => n3358);
   U401 : MUX2_X1 port map( A => n706, B => n1091, S => n1074, Z => n3357);
   U402 : MUX2_X1 port map( A => n707, B => n1092, S => n1074, Z => n3356);
   U403 : MUX2_X1 port map( A => n708, B => n1093, S => n1074, Z => n3355);
   U404 : MUX2_X1 port map( A => n709, B => n1094, S => n1074, Z => n3354);
   U405 : MUX2_X1 port map( A => n710, B => n1095, S => n1074, Z => n3353);
   U406 : MUX2_X1 port map( A => n711, B => n1096, S => n1074, Z => n3352);
   U407 : MUX2_X1 port map( A => n712, B => n1097, S => n1074, Z => n3351);
   U408 : MUX2_X1 port map( A => n713, B => n1098, S => n1074, Z => n3350);
   U409 : MUX2_X1 port map( A => n714, B => n1099, S => n1074, Z => n3349);
   U410 : MUX2_X1 port map( A => n715, B => n1100, S => n1074, Z => n3348);
   U411 : MUX2_X1 port map( A => n716, B => n1101, S => n1074, Z => n3347);
   U412 : MUX2_X1 port map( A => n717, B => n1102, S => n1074, Z => n3346);
   U413 : MUX2_X1 port map( A => n718, B => n1103, S => n1074, Z => n3345);
   U414 : MUX2_X1 port map( A => n719, B => n1104, S => n1074, Z => n3344);
   U415 : MUX2_X1 port map( A => n720, B => n1105, S => n1074, Z => n3343);
   U416 : MUX2_X1 port map( A => n721, B => n1106, S => n1074, Z => n3342);
   U417 : MUX2_X1 port map( A => n722, B => n1107, S => n1074, Z => n3341);
   U418 : MUX2_X1 port map( A => n723, B => n1108, S => n1074, Z => n3340);
   U419 : MUX2_X1 port map( A => n724, B => n1109, S => n1074, Z => n3339);
   U420 : MUX2_X1 port map( A => n725, B => n1110, S => n1074, Z => n3338);
   U421 : MUX2_X1 port map( A => n726, B => n1111, S => n1074, Z => n3337);
   U422 : MUX2_X1 port map( A => n727, B => n1112, S => n1074, Z => n3336);
   U423 : MUX2_X1 port map( A => n728, B => n1113, S => n1074, Z => n3335);
   U424 : MUX2_X1 port map( A => n729, B => n1114, S => n1074, Z => n3334);
   U425 : MUX2_X1 port map( A => n730, B => n1115, S => n1074, Z => n3333);
   U426 : MUX2_X1 port map( A => n731, B => n1116, S => n1074, Z => n3332);
   U427 : MUX2_X1 port map( A => n732, B => n1117, S => n1074, Z => n3331);
   U428 : MUX2_X1 port map( A => n733, B => n1118, S => n1074, Z => n3330);
   U429 : MUX2_X1 port map( A => n734, B => n1119, S => n1074, Z => n3329);
   U430 : MUX2_X1 port map( A => n735, B => n1120, S => n1074, Z => n3328);
   U431 : MUX2_X1 port map( A => n736, B => n1121, S => n1074, Z => n3327);
   U432 : OAI21_X1 port map( B1 => n1123, B2 => n1141, A => RST, ZN => n1140);
   U433 : MUX2_X1 port map( A => n321, B => n1089, S => n1068, Z => n3326);
   U434 : MUX2_X1 port map( A => n322, B => n1091, S => n1068, Z => n3325);
   U435 : MUX2_X1 port map( A => n323, B => n1092, S => n1068, Z => n3324);
   U436 : MUX2_X1 port map( A => n324, B => n1093, S => n1068, Z => n3323);
   U437 : MUX2_X1 port map( A => n325, B => n1094, S => n1068, Z => n3322);
   U438 : MUX2_X1 port map( A => n326, B => n1095, S => n1068, Z => n3321);
   U439 : MUX2_X1 port map( A => n327, B => n1096, S => n1068, Z => n3320);
   U440 : MUX2_X1 port map( A => n328, B => n1097, S => n1068, Z => n3319);
   U441 : MUX2_X1 port map( A => n329, B => n1098, S => n1068, Z => n3318);
   U442 : MUX2_X1 port map( A => n330, B => n1099, S => n1068, Z => n3317);
   U443 : MUX2_X1 port map( A => n331, B => n1100, S => n1068, Z => n3316);
   U444 : MUX2_X1 port map( A => n332, B => n1101, S => n1068, Z => n3315);
   U445 : MUX2_X1 port map( A => n333, B => n1102, S => n1068, Z => n3314);
   U446 : MUX2_X1 port map( A => n334, B => n1103, S => n1068, Z => n3313);
   U447 : MUX2_X1 port map( A => n335, B => n1104, S => n1068, Z => n3312);
   U448 : MUX2_X1 port map( A => n336, B => n1105, S => n1068, Z => n3311);
   U449 : MUX2_X1 port map( A => n337, B => n1106, S => n1068, Z => n3310);
   U450 : MUX2_X1 port map( A => n338, B => n1107, S => n1068, Z => n3309);
   U451 : MUX2_X1 port map( A => n339, B => n1108, S => n1068, Z => n3308);
   U452 : MUX2_X1 port map( A => n340, B => n1109, S => n1068, Z => n3307);
   U453 : MUX2_X1 port map( A => n341, B => n1110, S => n1068, Z => n3306);
   U454 : MUX2_X1 port map( A => n342, B => n1111, S => n1068, Z => n3305);
   U455 : MUX2_X1 port map( A => n343, B => n1112, S => n1068, Z => n3304);
   U456 : MUX2_X1 port map( A => n344, B => n1113, S => n1068, Z => n3303);
   U457 : MUX2_X1 port map( A => n345, B => n1114, S => n1068, Z => n3302);
   U458 : MUX2_X1 port map( A => n346, B => n1115, S => n1068, Z => n3301);
   U459 : MUX2_X1 port map( A => n347, B => n1116, S => n1068, Z => n3300);
   U460 : MUX2_X1 port map( A => n348, B => n1117, S => n1068, Z => n3299);
   U461 : MUX2_X1 port map( A => n349, B => n1118, S => n1068, Z => n3298);
   U462 : MUX2_X1 port map( A => n350, B => n1119, S => n1068, Z => n3297);
   U463 : MUX2_X1 port map( A => n351, B => n1120, S => n1068, Z => n3296);
   U464 : MUX2_X1 port map( A => n352, B => n1121, S => n1068, Z => n3295);
   U465 : OAI21_X1 port map( B1 => n1125, B2 => n1141, A => RST, ZN => n1142);
   U466 : MUX2_X1 port map( A => n4020, B => n1089, S => n1070, Z => n3294);
   U467 : MUX2_X1 port map( A => n4019, B => n1091, S => n1070, Z => n3293);
   U468 : MUX2_X1 port map( A => n4018, B => n1092, S => n1070, Z => n3292);
   U469 : MUX2_X1 port map( A => n4017, B => n1093, S => n1070, Z => n3291);
   U470 : MUX2_X1 port map( A => n4016, B => n1094, S => n1070, Z => n3290);
   U471 : MUX2_X1 port map( A => n4015, B => n1095, S => n1070, Z => n3289);
   U472 : MUX2_X1 port map( A => n4014, B => n1096, S => n1070, Z => n3288);
   U473 : MUX2_X1 port map( A => n4013, B => n1097, S => n1070, Z => n3287);
   U474 : MUX2_X1 port map( A => n4012, B => n1098, S => n1070, Z => n3286);
   U475 : MUX2_X1 port map( A => n4011, B => n1099, S => n1070, Z => n3285);
   U476 : MUX2_X1 port map( A => n4010, B => n1100, S => n1070, Z => n3284);
   U477 : MUX2_X1 port map( A => n4009, B => n1101, S => n1070, Z => n3283);
   U478 : MUX2_X1 port map( A => n4008, B => n1102, S => n1070, Z => n3282);
   U479 : MUX2_X1 port map( A => n4007, B => n1103, S => n1070, Z => n3281);
   U480 : MUX2_X1 port map( A => n4006, B => n1104, S => n1070, Z => n3280);
   U481 : MUX2_X1 port map( A => n4005, B => n1105, S => n1070, Z => n3279);
   U482 : MUX2_X1 port map( A => n4004, B => n1106, S => n1070, Z => n3278);
   U483 : MUX2_X1 port map( A => n4003, B => n1107, S => n1070, Z => n3277);
   U484 : MUX2_X1 port map( A => n4002, B => n1108, S => n1070, Z => n3276);
   U485 : MUX2_X1 port map( A => n4001, B => n1109, S => n1070, Z => n3275);
   U486 : MUX2_X1 port map( A => n4000, B => n1110, S => n1070, Z => n3274);
   U487 : MUX2_X1 port map( A => n3999, B => n1111, S => n1070, Z => n3273);
   U488 : MUX2_X1 port map( A => n3998, B => n1112, S => n1070, Z => n3272);
   U489 : MUX2_X1 port map( A => n3997, B => n1113, S => n1070, Z => n3271);
   U490 : MUX2_X1 port map( A => n3996, B => n1114, S => n1070, Z => n3270);
   U491 : MUX2_X1 port map( A => n3995, B => n1115, S => n1070, Z => n3269);
   U492 : MUX2_X1 port map( A => n3994, B => n1116, S => n1070, Z => n3268);
   U493 : MUX2_X1 port map( A => n3993, B => n1117, S => n1070, Z => n3267);
   U494 : MUX2_X1 port map( A => n3992, B => n1118, S => n1070, Z => n3266);
   U495 : MUX2_X1 port map( A => n3991, B => n1119, S => n1070, Z => n3265);
   U496 : MUX2_X1 port map( A => n3990, B => n1120, S => n1070, Z => n3264);
   U497 : MUX2_X1 port map( A => n3989, B => n1121, S => n1070, Z => n3263);
   U498 : OAI21_X1 port map( B1 => n1127, B2 => n1141, A => RST, ZN => n1143);
   U499 : MUX2_X1 port map( A => n3988, B => n1089, S => n1064, Z => n3262);
   U500 : MUX2_X1 port map( A => n3987, B => n1091, S => n1064, Z => n3261);
   U501 : MUX2_X1 port map( A => n3986, B => n1092, S => n1064, Z => n3260);
   U502 : MUX2_X1 port map( A => n3985, B => n1093, S => n1064, Z => n3259);
   U503 : MUX2_X1 port map( A => n3984, B => n1094, S => n1064, Z => n3258);
   U504 : MUX2_X1 port map( A => n3983, B => n1095, S => n1064, Z => n3257);
   U505 : MUX2_X1 port map( A => n3982, B => n1096, S => n1064, Z => n3256);
   U506 : MUX2_X1 port map( A => n3981, B => n1097, S => n1064, Z => n3255);
   U507 : MUX2_X1 port map( A => n3980, B => n1098, S => n1064, Z => n3254);
   U508 : MUX2_X1 port map( A => n3979, B => n1099, S => n1064, Z => n3253);
   U509 : MUX2_X1 port map( A => n3978, B => n1100, S => n1064, Z => n3252);
   U510 : MUX2_X1 port map( A => n3977, B => n1101, S => n1064, Z => n3251);
   U511 : MUX2_X1 port map( A => n3976, B => n1102, S => n1064, Z => n3250);
   U512 : MUX2_X1 port map( A => n3975, B => n1103, S => n1064, Z => n3249);
   U513 : MUX2_X1 port map( A => n3974, B => n1104, S => n1064, Z => n3248);
   U514 : MUX2_X1 port map( A => n3973, B => n1105, S => n1064, Z => n3247);
   U515 : MUX2_X1 port map( A => n3972, B => n1106, S => n1064, Z => n3246);
   U516 : MUX2_X1 port map( A => n3971, B => n1107, S => n1064, Z => n3245);
   U517 : MUX2_X1 port map( A => n3970, B => n1108, S => n1064, Z => n3244);
   U518 : MUX2_X1 port map( A => n3969, B => n1109, S => n1064, Z => n3243);
   U519 : MUX2_X1 port map( A => n3968, B => n1110, S => n1064, Z => n3242);
   U520 : MUX2_X1 port map( A => n3967, B => n1111, S => n1064, Z => n3241);
   U521 : MUX2_X1 port map( A => n3966, B => n1112, S => n1064, Z => n3240);
   U522 : MUX2_X1 port map( A => n3965, B => n1113, S => n1064, Z => n3239);
   U523 : MUX2_X1 port map( A => n3964, B => n1114, S => n1064, Z => n3238);
   U524 : MUX2_X1 port map( A => n3963, B => n1115, S => n1064, Z => n3237);
   U525 : MUX2_X1 port map( A => n3962, B => n1116, S => n1064, Z => n3236);
   U526 : MUX2_X1 port map( A => n3961, B => n1117, S => n1064, Z => n3235);
   U527 : MUX2_X1 port map( A => n3960, B => n1118, S => n1064, Z => n3234);
   U528 : MUX2_X1 port map( A => n3959, B => n1119, S => n1064, Z => n3233);
   U529 : MUX2_X1 port map( A => n3958, B => n1120, S => n1064, Z => n3232);
   U530 : MUX2_X1 port map( A => n3957, B => n1121, S => n1064, Z => n3231);
   U531 : OAI21_X1 port map( B1 => n1129, B2 => n1141, A => RST, ZN => n1144);
   U532 : MUX2_X1 port map( A => n737, B => n1089, S => n1066, Z => n3230);
   U533 : MUX2_X1 port map( A => n738, B => n1091, S => n1066, Z => n3229);
   U534 : MUX2_X1 port map( A => n739, B => n1092, S => n1066, Z => n3228);
   U535 : MUX2_X1 port map( A => n740, B => n1093, S => n1066, Z => n3227);
   U536 : MUX2_X1 port map( A => n741, B => n1094, S => n1066, Z => n3226);
   U537 : MUX2_X1 port map( A => n742, B => n1095, S => n1066, Z => n3225);
   U538 : MUX2_X1 port map( A => n743, B => n1096, S => n1066, Z => n3224);
   U539 : MUX2_X1 port map( A => n744, B => n1097, S => n1066, Z => n3223);
   U540 : MUX2_X1 port map( A => n745, B => n1098, S => n1066, Z => n3222);
   U541 : MUX2_X1 port map( A => n746, B => n1099, S => n1066, Z => n3221);
   U542 : MUX2_X1 port map( A => n747, B => n1100, S => n1066, Z => n3220);
   U543 : MUX2_X1 port map( A => n748, B => n1101, S => n1066, Z => n3219);
   U544 : MUX2_X1 port map( A => n749, B => n1102, S => n1066, Z => n3218);
   U545 : MUX2_X1 port map( A => n750, B => n1103, S => n1066, Z => n3217);
   U546 : MUX2_X1 port map( A => n751, B => n1104, S => n1066, Z => n3216);
   U547 : MUX2_X1 port map( A => n752, B => n1105, S => n1066, Z => n3215);
   U548 : MUX2_X1 port map( A => n753, B => n1106, S => n1066, Z => n3214);
   U549 : MUX2_X1 port map( A => n754, B => n1107, S => n1066, Z => n3213);
   U550 : MUX2_X1 port map( A => n755, B => n1108, S => n1066, Z => n3212);
   U551 : MUX2_X1 port map( A => n756, B => n1109, S => n1066, Z => n3211);
   U552 : MUX2_X1 port map( A => n757, B => n1110, S => n1066, Z => n3210);
   U553 : MUX2_X1 port map( A => n758, B => n1111, S => n1066, Z => n3209);
   U554 : MUX2_X1 port map( A => n759, B => n1112, S => n1066, Z => n3208);
   U555 : MUX2_X1 port map( A => n760, B => n1113, S => n1066, Z => n3207);
   U556 : MUX2_X1 port map( A => n761, B => n1114, S => n1066, Z => n3206);
   U557 : MUX2_X1 port map( A => n762, B => n1115, S => n1066, Z => n3205);
   U558 : MUX2_X1 port map( A => n763, B => n1116, S => n1066, Z => n3204);
   U559 : MUX2_X1 port map( A => n764, B => n1117, S => n1066, Z => n3203);
   U560 : MUX2_X1 port map( A => n765, B => n1118, S => n1066, Z => n3202);
   U561 : MUX2_X1 port map( A => n766, B => n1119, S => n1066, Z => n3201);
   U562 : MUX2_X1 port map( A => n767, B => n1120, S => n1066, Z => n3200);
   U563 : MUX2_X1 port map( A => n768, B => n1121, S => n1066, Z => n3199);
   U564 : OAI21_X1 port map( B1 => n1131, B2 => n1141, A => RST, ZN => n1145);
   U565 : MUX2_X1 port map( A => n353, B => n1089, S => n1060, Z => n3198);
   U566 : MUX2_X1 port map( A => n354, B => n1091, S => n1060, Z => n3197);
   U567 : MUX2_X1 port map( A => n355, B => n1092, S => n1060, Z => n3196);
   U568 : MUX2_X1 port map( A => n356, B => n1093, S => n1060, Z => n3195);
   U569 : MUX2_X1 port map( A => n357, B => n1094, S => n1060, Z => n3194);
   U570 : MUX2_X1 port map( A => n358, B => n1095, S => n1060, Z => n3193);
   U571 : MUX2_X1 port map( A => n359, B => n1096, S => n1060, Z => n3192);
   U572 : MUX2_X1 port map( A => n360, B => n1097, S => n1060, Z => n3191);
   U573 : MUX2_X1 port map( A => n361, B => n1098, S => n1060, Z => n3190);
   U574 : MUX2_X1 port map( A => n362, B => n1099, S => n1060, Z => n3189);
   U575 : MUX2_X1 port map( A => n363, B => n1100, S => n1060, Z => n3188);
   U576 : MUX2_X1 port map( A => n364, B => n1101, S => n1060, Z => n3187);
   U577 : MUX2_X1 port map( A => n365, B => n1102, S => n1060, Z => n3186);
   U578 : MUX2_X1 port map( A => n366, B => n1103, S => n1060, Z => n3185);
   U579 : MUX2_X1 port map( A => n367, B => n1104, S => n1060, Z => n3184);
   U580 : MUX2_X1 port map( A => n368, B => n1105, S => n1060, Z => n3183);
   U581 : MUX2_X1 port map( A => n369, B => n1106, S => n1060, Z => n3182);
   U582 : MUX2_X1 port map( A => n370, B => n1107, S => n1060, Z => n3181);
   U583 : MUX2_X1 port map( A => n371, B => n1108, S => n1060, Z => n3180);
   U584 : MUX2_X1 port map( A => n372, B => n1109, S => n1060, Z => n3179);
   U585 : MUX2_X1 port map( A => n373, B => n1110, S => n1060, Z => n3178);
   U586 : MUX2_X1 port map( A => n374, B => n1111, S => n1060, Z => n3177);
   U587 : MUX2_X1 port map( A => n375, B => n1112, S => n1060, Z => n3176);
   U588 : MUX2_X1 port map( A => n376, B => n1113, S => n1060, Z => n3175);
   U589 : MUX2_X1 port map( A => n377, B => n1114, S => n1060, Z => n3174);
   U590 : MUX2_X1 port map( A => n378, B => n1115, S => n1060, Z => n3173);
   U591 : MUX2_X1 port map( A => n379, B => n1116, S => n1060, Z => n3172);
   U592 : MUX2_X1 port map( A => n380, B => n1117, S => n1060, Z => n3171);
   U593 : MUX2_X1 port map( A => n381, B => n1118, S => n1060, Z => n3170);
   U594 : MUX2_X1 port map( A => n382, B => n1119, S => n1060, Z => n3169);
   U595 : MUX2_X1 port map( A => n383, B => n1120, S => n1060, Z => n3168);
   U596 : MUX2_X1 port map( A => n384, B => n1121, S => n1060, Z => n3167);
   U597 : OAI21_X1 port map( B1 => n1133, B2 => n1141, A => RST, ZN => n1146);
   U598 : MUX2_X1 port map( A => n3956, B => n1089, S => n1062, Z => n3166);
   U599 : MUX2_X1 port map( A => n3955, B => n1091, S => n1062, Z => n3165);
   U600 : MUX2_X1 port map( A => n3954, B => n1092, S => n1062, Z => n3164);
   U601 : MUX2_X1 port map( A => n3953, B => n1093, S => n1062, Z => n3163);
   U602 : MUX2_X1 port map( A => n3952, B => n1094, S => n1062, Z => n3162);
   U603 : MUX2_X1 port map( A => n3951, B => n1095, S => n1062, Z => n3161);
   U604 : MUX2_X1 port map( A => n3950, B => n1096, S => n1062, Z => n3160);
   U605 : MUX2_X1 port map( A => n3949, B => n1097, S => n1062, Z => n3159);
   U606 : MUX2_X1 port map( A => n3948, B => n1098, S => n1062, Z => n3158);
   U607 : MUX2_X1 port map( A => n3947, B => n1099, S => n1062, Z => n3157);
   U608 : MUX2_X1 port map( A => n3946, B => n1100, S => n1062, Z => n3156);
   U609 : MUX2_X1 port map( A => n3945, B => n1101, S => n1062, Z => n3155);
   U610 : MUX2_X1 port map( A => n3944, B => n1102, S => n1062, Z => n3154);
   U611 : MUX2_X1 port map( A => n3943, B => n1103, S => n1062, Z => n3153);
   U612 : MUX2_X1 port map( A => n3942, B => n1104, S => n1062, Z => n3152);
   U613 : MUX2_X1 port map( A => n3941, B => n1105, S => n1062, Z => n3151);
   U614 : MUX2_X1 port map( A => n3940, B => n1106, S => n1062, Z => n3150);
   U615 : MUX2_X1 port map( A => n3939, B => n1107, S => n1062, Z => n3149);
   U616 : MUX2_X1 port map( A => n3938, B => n1108, S => n1062, Z => n3148);
   U617 : MUX2_X1 port map( A => n3937, B => n1109, S => n1062, Z => n3147);
   U618 : MUX2_X1 port map( A => n3936, B => n1110, S => n1062, Z => n3146);
   U619 : MUX2_X1 port map( A => n3935, B => n1111, S => n1062, Z => n3145);
   U620 : MUX2_X1 port map( A => n3934, B => n1112, S => n1062, Z => n3144);
   U621 : MUX2_X1 port map( A => n3933, B => n1113, S => n1062, Z => n3143);
   U622 : MUX2_X1 port map( A => n3932, B => n1114, S => n1062, Z => n3142);
   U623 : MUX2_X1 port map( A => n3931, B => n1115, S => n1062, Z => n3141);
   U624 : MUX2_X1 port map( A => n3930, B => n1116, S => n1062, Z => n3140);
   U625 : MUX2_X1 port map( A => n3929, B => n1117, S => n1062, Z => n3139);
   U626 : MUX2_X1 port map( A => n3928, B => n1118, S => n1062, Z => n3138);
   U627 : MUX2_X1 port map( A => n3927, B => n1119, S => n1062, Z => n3137);
   U628 : MUX2_X1 port map( A => n3926, B => n1120, S => n1062, Z => n3136);
   U629 : MUX2_X1 port map( A => n3925, B => n1121, S => n1062, Z => n3135);
   U630 : OAI21_X1 port map( B1 => n1135, B2 => n1141, A => RST, ZN => n1147);
   U631 : MUX2_X1 port map( A => n3924, B => n1089, S => n1056, Z => n3134);
   U632 : MUX2_X1 port map( A => n3923, B => n1091, S => n1056, Z => n3133);
   U633 : MUX2_X1 port map( A => n3922, B => n1092, S => n1056, Z => n3132);
   U634 : MUX2_X1 port map( A => n3921, B => n1093, S => n1056, Z => n3131);
   U635 : MUX2_X1 port map( A => n3920, B => n1094, S => n1056, Z => n3130);
   U636 : MUX2_X1 port map( A => n3919, B => n1095, S => n1056, Z => n3129);
   U637 : MUX2_X1 port map( A => n3918, B => n1096, S => n1056, Z => n3128);
   U638 : MUX2_X1 port map( A => n3917, B => n1097, S => n1056, Z => n3127);
   U639 : MUX2_X1 port map( A => n3916, B => n1098, S => n1056, Z => n3126);
   U640 : MUX2_X1 port map( A => n3915, B => n1099, S => n1056, Z => n3125);
   U641 : MUX2_X1 port map( A => n3914, B => n1100, S => n1056, Z => n3124);
   U642 : MUX2_X1 port map( A => n3913, B => n1101, S => n1056, Z => n3123);
   U643 : MUX2_X1 port map( A => n3912, B => n1102, S => n1056, Z => n3122);
   U644 : MUX2_X1 port map( A => n3911, B => n1103, S => n1056, Z => n3121);
   U645 : MUX2_X1 port map( A => n3910, B => n1104, S => n1056, Z => n3120);
   U646 : MUX2_X1 port map( A => n3909, B => n1105, S => n1056, Z => n3119);
   U647 : MUX2_X1 port map( A => n3908, B => n1106, S => n1056, Z => n3118);
   U648 : MUX2_X1 port map( A => n3907, B => n1107, S => n1056, Z => n3117);
   U649 : MUX2_X1 port map( A => n3906, B => n1108, S => n1056, Z => n3116);
   U650 : MUX2_X1 port map( A => n3905, B => n1109, S => n1056, Z => n3115);
   U651 : MUX2_X1 port map( A => n3904, B => n1110, S => n1056, Z => n3114);
   U652 : MUX2_X1 port map( A => n3903, B => n1111, S => n1056, Z => n3113);
   U653 : MUX2_X1 port map( A => n3902, B => n1112, S => n1056, Z => n3112);
   U654 : MUX2_X1 port map( A => n3901, B => n1113, S => n1056, Z => n3111);
   U655 : MUX2_X1 port map( A => n3900, B => n1114, S => n1056, Z => n3110);
   U656 : MUX2_X1 port map( A => n3899, B => n1115, S => n1056, Z => n3109);
   U657 : MUX2_X1 port map( A => n3898, B => n1116, S => n1056, Z => n3108);
   U658 : MUX2_X1 port map( A => n3897, B => n1117, S => n1056, Z => n3107);
   U659 : MUX2_X1 port map( A => n3896, B => n1118, S => n1056, Z => n3106);
   U660 : MUX2_X1 port map( A => n3895, B => n1119, S => n1056, Z => n3105);
   U661 : MUX2_X1 port map( A => n3894, B => n1120, S => n1056, Z => n3104);
   U662 : MUX2_X1 port map( A => n3893, B => n1121, S => n1056, Z => n3103);
   U663 : OAI21_X1 port map( B1 => n1137, B2 => n1141, A => RST, ZN => n1148);
   U664 : NAND3_X1 port map( A1 => WR, A2 => n1139, A3 => ADD_WR(3), ZN => 
                           n1141);
   U665 : INV_X1 port map( A => ADD_WR(4), ZN => n1139);
   U666 : MUX2_X1 port map( A => n769, B => n1089, S => n1058, Z => n3102);
   U667 : MUX2_X1 port map( A => n770, B => n1091, S => n1058, Z => n3101);
   U668 : MUX2_X1 port map( A => n771, B => n1092, S => n1058, Z => n3100);
   U669 : MUX2_X1 port map( A => n772, B => n1093, S => n1058, Z => n3099);
   U670 : MUX2_X1 port map( A => n773, B => n1094, S => n1058, Z => n3098);
   U671 : MUX2_X1 port map( A => n774, B => n1095, S => n1058, Z => n3097);
   U672 : MUX2_X1 port map( A => n775, B => n1096, S => n1058, Z => n3096);
   U673 : MUX2_X1 port map( A => n776, B => n1097, S => n1058, Z => n3095);
   U674 : MUX2_X1 port map( A => n777, B => n1098, S => n1058, Z => n3094);
   U675 : MUX2_X1 port map( A => n778, B => n1099, S => n1058, Z => n3093);
   U676 : MUX2_X1 port map( A => n779, B => n1100, S => n1058, Z => n3092);
   U677 : MUX2_X1 port map( A => n780, B => n1101, S => n1058, Z => n3091);
   U678 : MUX2_X1 port map( A => n781, B => n1102, S => n1058, Z => n3090);
   U679 : MUX2_X1 port map( A => n782, B => n1103, S => n1058, Z => n3089);
   U680 : MUX2_X1 port map( A => n783, B => n1104, S => n1058, Z => n3088);
   U681 : MUX2_X1 port map( A => n784, B => n1105, S => n1058, Z => n3087);
   U682 : MUX2_X1 port map( A => n785, B => n1106, S => n1058, Z => n3086);
   U683 : MUX2_X1 port map( A => n786, B => n1107, S => n1058, Z => n3085);
   U684 : MUX2_X1 port map( A => n787, B => n1108, S => n1058, Z => n3084);
   U685 : MUX2_X1 port map( A => n788, B => n1109, S => n1058, Z => n3083);
   U686 : MUX2_X1 port map( A => n789, B => n1110, S => n1058, Z => n3082);
   U687 : MUX2_X1 port map( A => n790, B => n1111, S => n1058, Z => n3081);
   U688 : MUX2_X1 port map( A => n791, B => n1112, S => n1058, Z => n3080);
   U689 : MUX2_X1 port map( A => n792, B => n1113, S => n1058, Z => n3079);
   U690 : MUX2_X1 port map( A => n793, B => n1114, S => n1058, Z => n3078);
   U691 : MUX2_X1 port map( A => n794, B => n1115, S => n1058, Z => n3077);
   U692 : MUX2_X1 port map( A => n795, B => n1116, S => n1058, Z => n3076);
   U693 : MUX2_X1 port map( A => n796, B => n1117, S => n1058, Z => n3075);
   U694 : MUX2_X1 port map( A => n797, B => n1118, S => n1058, Z => n3074);
   U695 : MUX2_X1 port map( A => n798, B => n1119, S => n1058, Z => n3073);
   U696 : MUX2_X1 port map( A => n799, B => n1120, S => n1058, Z => n3072);
   U697 : MUX2_X1 port map( A => n800, B => n1121, S => n1058, Z => n3071);
   U698 : OAI21_X1 port map( B1 => n1123, B2 => n1150, A => RST, ZN => n1149);
   U699 : MUX2_X1 port map( A => n449, B => n1089, S => n1052, Z => n3070);
   U700 : MUX2_X1 port map( A => n450, B => n1091, S => n1052, Z => n3069);
   U701 : MUX2_X1 port map( A => n451, B => n1092, S => n1052, Z => n3068);
   U702 : MUX2_X1 port map( A => n452, B => n1093, S => n1052, Z => n3067);
   U703 : MUX2_X1 port map( A => n453, B => n1094, S => n1052, Z => n3066);
   U704 : MUX2_X1 port map( A => n454, B => n1095, S => n1052, Z => n3065);
   U705 : MUX2_X1 port map( A => n455, B => n1096, S => n1052, Z => n3064);
   U706 : MUX2_X1 port map( A => n456, B => n1097, S => n1052, Z => n3063);
   U707 : MUX2_X1 port map( A => n457, B => n1098, S => n1052, Z => n3062);
   U708 : MUX2_X1 port map( A => n458, B => n1099, S => n1052, Z => n3061);
   U709 : MUX2_X1 port map( A => n459, B => n1100, S => n1052, Z => n3060);
   U710 : MUX2_X1 port map( A => n460, B => n1101, S => n1052, Z => n3059);
   U711 : MUX2_X1 port map( A => n461, B => n1102, S => n1052, Z => n3058);
   U712 : MUX2_X1 port map( A => n462, B => n1103, S => n1052, Z => n3057);
   U713 : MUX2_X1 port map( A => n463, B => n1104, S => n1052, Z => n3056);
   U714 : MUX2_X1 port map( A => n464, B => n1105, S => n1052, Z => n3055);
   U715 : MUX2_X1 port map( A => n465, B => n1106, S => n1052, Z => n3054);
   U716 : MUX2_X1 port map( A => n466, B => n1107, S => n1052, Z => n3053);
   U717 : MUX2_X1 port map( A => n467, B => n1108, S => n1052, Z => n3052);
   U718 : MUX2_X1 port map( A => n468, B => n1109, S => n1052, Z => n3051);
   U719 : MUX2_X1 port map( A => n469, B => n1110, S => n1052, Z => n3050);
   U720 : MUX2_X1 port map( A => n470, B => n1111, S => n1052, Z => n3049);
   U721 : MUX2_X1 port map( A => n471, B => n1112, S => n1052, Z => n3048);
   U722 : MUX2_X1 port map( A => n472, B => n1113, S => n1052, Z => n3047);
   U723 : MUX2_X1 port map( A => n473, B => n1114, S => n1052, Z => n3046);
   U724 : MUX2_X1 port map( A => n474, B => n1115, S => n1052, Z => n3045);
   U725 : MUX2_X1 port map( A => n475, B => n1116, S => n1052, Z => n3044);
   U726 : MUX2_X1 port map( A => n476, B => n1117, S => n1052, Z => n3043);
   U727 : MUX2_X1 port map( A => n477, B => n1118, S => n1052, Z => n3042);
   U728 : MUX2_X1 port map( A => n478, B => n1119, S => n1052, Z => n3041);
   U729 : MUX2_X1 port map( A => n479, B => n1120, S => n1052, Z => n3040);
   U730 : MUX2_X1 port map( A => n480, B => n1121, S => n1052, Z => n3039);
   U731 : OAI21_X1 port map( B1 => n1125, B2 => n1150, A => RST, ZN => n1151);
   U732 : MUX2_X1 port map( A => n3892, B => n1089, S => n1054, Z => n3038);
   U733 : MUX2_X1 port map( A => n3891, B => n1091, S => n1054, Z => n3037);
   U734 : MUX2_X1 port map( A => n3890, B => n1092, S => n1054, Z => n3036);
   U735 : MUX2_X1 port map( A => n3889, B => n1093, S => n1054, Z => n3035);
   U736 : MUX2_X1 port map( A => n3888, B => n1094, S => n1054, Z => n3034);
   U737 : MUX2_X1 port map( A => n3887, B => n1095, S => n1054, Z => n3033);
   U738 : MUX2_X1 port map( A => n3886, B => n1096, S => n1054, Z => n3032);
   U739 : MUX2_X1 port map( A => n3885, B => n1097, S => n1054, Z => n3031);
   U740 : MUX2_X1 port map( A => n3884, B => n1098, S => n1054, Z => n3030);
   U741 : MUX2_X1 port map( A => n3883, B => n1099, S => n1054, Z => n3029);
   U742 : MUX2_X1 port map( A => n3882, B => n1100, S => n1054, Z => n3028);
   U743 : MUX2_X1 port map( A => n3881, B => n1101, S => n1054, Z => n3027);
   U744 : MUX2_X1 port map( A => n3880, B => n1102, S => n1054, Z => n3026);
   U745 : MUX2_X1 port map( A => n3879, B => n1103, S => n1054, Z => n3025);
   U746 : MUX2_X1 port map( A => n3878, B => n1104, S => n1054, Z => n3024);
   U747 : MUX2_X1 port map( A => n3877, B => n1105, S => n1054, Z => n3023);
   U748 : MUX2_X1 port map( A => n3876, B => n1106, S => n1054, Z => n3022);
   U749 : MUX2_X1 port map( A => n3875, B => n1107, S => n1054, Z => n3021);
   U750 : MUX2_X1 port map( A => n3874, B => n1108, S => n1054, Z => n3020);
   U751 : MUX2_X1 port map( A => n3873, B => n1109, S => n1054, Z => n3019);
   U752 : MUX2_X1 port map( A => n3872, B => n1110, S => n1054, Z => n3018);
   U753 : MUX2_X1 port map( A => n3871, B => n1111, S => n1054, Z => n3017);
   U754 : MUX2_X1 port map( A => n3870, B => n1112, S => n1054, Z => n3016);
   U755 : MUX2_X1 port map( A => n3869, B => n1113, S => n1054, Z => n3015);
   U756 : MUX2_X1 port map( A => n3868, B => n1114, S => n1054, Z => n3014);
   U757 : MUX2_X1 port map( A => n3867, B => n1115, S => n1054, Z => n3013);
   U758 : MUX2_X1 port map( A => n3866, B => n1116, S => n1054, Z => n3012);
   U759 : MUX2_X1 port map( A => n3865, B => n1117, S => n1054, Z => n3011);
   U760 : MUX2_X1 port map( A => n3864, B => n1118, S => n1054, Z => n3010);
   U761 : MUX2_X1 port map( A => n3863, B => n1119, S => n1054, Z => n3009);
   U762 : MUX2_X1 port map( A => n3862, B => n1120, S => n1054, Z => n3008);
   U763 : MUX2_X1 port map( A => n3861, B => n1121, S => n1054, Z => n3007);
   U764 : OAI21_X1 port map( B1 => n1127, B2 => n1150, A => RST, ZN => n1152);
   U765 : MUX2_X1 port map( A => n3860, B => n1089, S => n1026, Z => n3006);
   U766 : MUX2_X1 port map( A => n3859, B => n1091, S => n1026, Z => n3005);
   U767 : MUX2_X1 port map( A => n3858, B => n1092, S => n1026, Z => n3004);
   U768 : MUX2_X1 port map( A => n3857, B => n1093, S => n1026, Z => n3003);
   U769 : MUX2_X1 port map( A => n3856, B => n1094, S => n1026, Z => n3002);
   U770 : MUX2_X1 port map( A => n3855, B => n1095, S => n1026, Z => n3001);
   U771 : MUX2_X1 port map( A => n3854, B => n1096, S => n1026, Z => n3000);
   U772 : MUX2_X1 port map( A => n3853, B => n1097, S => n1026, Z => n2999);
   U773 : MUX2_X1 port map( A => n3852, B => n1098, S => n1026, Z => n2998);
   U774 : MUX2_X1 port map( A => n3851, B => n1099, S => n1026, Z => n2997);
   U775 : MUX2_X1 port map( A => n3850, B => n1100, S => n1026, Z => n2996);
   U776 : MUX2_X1 port map( A => n3849, B => n1101, S => n1026, Z => n2995);
   U777 : MUX2_X1 port map( A => n3848, B => n1102, S => n1026, Z => n2994);
   U778 : MUX2_X1 port map( A => n3847, B => n1103, S => n1026, Z => n2993);
   U779 : MUX2_X1 port map( A => n3846, B => n1104, S => n1026, Z => n2992);
   U780 : MUX2_X1 port map( A => n3845, B => n1105, S => n1026, Z => n2991);
   U781 : MUX2_X1 port map( A => n3844, B => n1106, S => n1026, Z => n2990);
   U782 : MUX2_X1 port map( A => n3843, B => n1107, S => n1026, Z => n2989);
   U783 : MUX2_X1 port map( A => n3842, B => n1108, S => n1026, Z => n2988);
   U784 : MUX2_X1 port map( A => n3841, B => n1109, S => n1026, Z => n2987);
   U785 : MUX2_X1 port map( A => n3840, B => n1110, S => n1026, Z => n2986);
   U786 : MUX2_X1 port map( A => n3839, B => n1111, S => n1026, Z => n2985);
   U787 : MUX2_X1 port map( A => n3838, B => n1112, S => n1026, Z => n2984);
   U788 : MUX2_X1 port map( A => n3837, B => n1113, S => n1026, Z => n2983);
   U789 : MUX2_X1 port map( A => n3836, B => n1114, S => n1026, Z => n2982);
   U790 : MUX2_X1 port map( A => n3835, B => n1115, S => n1026, Z => n2981);
   U791 : MUX2_X1 port map( A => n3834, B => n1116, S => n1026, Z => n2980);
   U792 : MUX2_X1 port map( A => n3833, B => n1117, S => n1026, Z => n2979);
   U793 : MUX2_X1 port map( A => n3832, B => n1118, S => n1026, Z => n2978);
   U794 : MUX2_X1 port map( A => n3831, B => n1119, S => n1026, Z => n2977);
   U795 : MUX2_X1 port map( A => n3830, B => n1120, S => n1026, Z => n2976);
   U796 : MUX2_X1 port map( A => n3829, B => n1121, S => n1026, Z => n2975);
   U797 : OAI21_X1 port map( B1 => n1129, B2 => n1150, A => RST, ZN => n1153);
   U798 : MUX2_X1 port map( A => n801, B => n1089, S => n1028, Z => n2974);
   U799 : MUX2_X1 port map( A => n802, B => n1091, S => n1028, Z => n2973);
   U800 : MUX2_X1 port map( A => n803, B => n1092, S => n1028, Z => n2972);
   U801 : MUX2_X1 port map( A => n804, B => n1093, S => n1028, Z => n2971);
   U802 : MUX2_X1 port map( A => n805, B => n1094, S => n1028, Z => n2970);
   U803 : MUX2_X1 port map( A => n806, B => n1095, S => n1028, Z => n2969);
   U804 : MUX2_X1 port map( A => n807, B => n1096, S => n1028, Z => n2968);
   U805 : MUX2_X1 port map( A => n808, B => n1097, S => n1028, Z => n2967);
   U806 : MUX2_X1 port map( A => n809, B => n1098, S => n1028, Z => n2966);
   U807 : MUX2_X1 port map( A => n810, B => n1099, S => n1028, Z => n2965);
   U808 : MUX2_X1 port map( A => n811, B => n1100, S => n1028, Z => n2964);
   U809 : MUX2_X1 port map( A => n812, B => n1101, S => n1028, Z => n2963);
   U810 : MUX2_X1 port map( A => n813, B => n1102, S => n1028, Z => n2962);
   U811 : MUX2_X1 port map( A => n814, B => n1103, S => n1028, Z => n2961);
   U812 : MUX2_X1 port map( A => n815, B => n1104, S => n1028, Z => n2960);
   U813 : MUX2_X1 port map( A => n816, B => n1105, S => n1028, Z => n2959);
   U814 : MUX2_X1 port map( A => n817, B => n1106, S => n1028, Z => n2958);
   U815 : MUX2_X1 port map( A => n818, B => n1107, S => n1028, Z => n2957);
   U816 : MUX2_X1 port map( A => n819, B => n1108, S => n1028, Z => n2956);
   U817 : MUX2_X1 port map( A => n820, B => n1109, S => n1028, Z => n2955);
   U818 : MUX2_X1 port map( A => n821, B => n1110, S => n1028, Z => n2954);
   U819 : MUX2_X1 port map( A => n822, B => n1111, S => n1028, Z => n2953);
   U820 : MUX2_X1 port map( A => n823, B => n1112, S => n1028, Z => n2952);
   U821 : MUX2_X1 port map( A => n824, B => n1113, S => n1028, Z => n2951);
   U822 : MUX2_X1 port map( A => n825, B => n1114, S => n1028, Z => n2950);
   U823 : MUX2_X1 port map( A => n826, B => n1115, S => n1028, Z => n2949);
   U824 : MUX2_X1 port map( A => n827, B => n1116, S => n1028, Z => n2948);
   U825 : MUX2_X1 port map( A => n828, B => n1117, S => n1028, Z => n2947);
   U826 : MUX2_X1 port map( A => n829, B => n1118, S => n1028, Z => n2946);
   U827 : MUX2_X1 port map( A => n830, B => n1119, S => n1028, Z => n2945);
   U828 : MUX2_X1 port map( A => n831, B => n1120, S => n1028, Z => n2944);
   U829 : MUX2_X1 port map( A => n832, B => n1121, S => n1028, Z => n2943);
   U830 : OAI21_X1 port map( B1 => n1131, B2 => n1150, A => RST, ZN => n1154);
   U831 : MUX2_X1 port map( A => n481, B => n1089, S => n1030, Z => n2942);
   U832 : MUX2_X1 port map( A => n482, B => n1091, S => n1030, Z => n2941);
   U833 : MUX2_X1 port map( A => n483, B => n1092, S => n1030, Z => n2940);
   U834 : MUX2_X1 port map( A => n484, B => n1093, S => n1030, Z => n2939);
   U835 : MUX2_X1 port map( A => n485, B => n1094, S => n1030, Z => n2938);
   U836 : MUX2_X1 port map( A => n486, B => n1095, S => n1030, Z => n2937);
   U837 : MUX2_X1 port map( A => n487, B => n1096, S => n1030, Z => n2936);
   U838 : MUX2_X1 port map( A => n488, B => n1097, S => n1030, Z => n2935);
   U839 : MUX2_X1 port map( A => n489, B => n1098, S => n1030, Z => n2934);
   U840 : MUX2_X1 port map( A => n490, B => n1099, S => n1030, Z => n2933);
   U841 : MUX2_X1 port map( A => n491, B => n1100, S => n1030, Z => n2932);
   U842 : MUX2_X1 port map( A => n492, B => n1101, S => n1030, Z => n2931);
   U843 : MUX2_X1 port map( A => n493, B => n1102, S => n1030, Z => n2930);
   U844 : MUX2_X1 port map( A => n494, B => n1103, S => n1030, Z => n2929);
   U845 : MUX2_X1 port map( A => n495, B => n1104, S => n1030, Z => n2928);
   U846 : MUX2_X1 port map( A => n496, B => n1105, S => n1030, Z => n2927);
   U847 : MUX2_X1 port map( A => n497, B => n1106, S => n1030, Z => n2926);
   U848 : MUX2_X1 port map( A => n498, B => n1107, S => n1030, Z => n2925);
   U849 : MUX2_X1 port map( A => n499, B => n1108, S => n1030, Z => n2924);
   U850 : MUX2_X1 port map( A => n500, B => n1109, S => n1030, Z => n2923);
   U851 : MUX2_X1 port map( A => n501, B => n1110, S => n1030, Z => n2922);
   U852 : MUX2_X1 port map( A => n502, B => n1111, S => n1030, Z => n2921);
   U853 : MUX2_X1 port map( A => n503, B => n1112, S => n1030, Z => n2920);
   U854 : MUX2_X1 port map( A => n504, B => n1113, S => n1030, Z => n2919);
   U855 : MUX2_X1 port map( A => n505, B => n1114, S => n1030, Z => n2918);
   U856 : MUX2_X1 port map( A => n506, B => n1115, S => n1030, Z => n2917);
   U857 : MUX2_X1 port map( A => n507, B => n1116, S => n1030, Z => n2916);
   U858 : MUX2_X1 port map( A => n508, B => n1117, S => n1030, Z => n2915);
   U859 : MUX2_X1 port map( A => n509, B => n1118, S => n1030, Z => n2914);
   U860 : MUX2_X1 port map( A => n510, B => n1119, S => n1030, Z => n2913);
   U861 : MUX2_X1 port map( A => n511, B => n1120, S => n1030, Z => n2912);
   U862 : MUX2_X1 port map( A => n512, B => n1121, S => n1030, Z => n2911);
   U863 : OAI21_X1 port map( B1 => n1133, B2 => n1150, A => RST, ZN => n1155);
   U864 : MUX2_X1 port map( A => n3828, B => n1089, S => n1032, Z => n2910);
   U865 : MUX2_X1 port map( A => n3827, B => n1091, S => n1032, Z => n2909);
   U866 : MUX2_X1 port map( A => n3826, B => n1092, S => n1032, Z => n2908);
   U867 : MUX2_X1 port map( A => n3825, B => n1093, S => n1032, Z => n2907);
   U868 : MUX2_X1 port map( A => n3824, B => n1094, S => n1032, Z => n2906);
   U869 : MUX2_X1 port map( A => n3823, B => n1095, S => n1032, Z => n2905);
   U870 : MUX2_X1 port map( A => n3822, B => n1096, S => n1032, Z => n2904);
   U871 : MUX2_X1 port map( A => n3821, B => n1097, S => n1032, Z => n2903);
   U872 : MUX2_X1 port map( A => n3820, B => n1098, S => n1032, Z => n2902);
   U873 : MUX2_X1 port map( A => n3819, B => n1099, S => n1032, Z => n2901);
   U874 : MUX2_X1 port map( A => n3818, B => n1100, S => n1032, Z => n2900);
   U875 : MUX2_X1 port map( A => n3817, B => n1101, S => n1032, Z => n2899);
   U876 : MUX2_X1 port map( A => n3816, B => n1102, S => n1032, Z => n2898);
   U877 : MUX2_X1 port map( A => n3815, B => n1103, S => n1032, Z => n2897);
   U878 : MUX2_X1 port map( A => n3814, B => n1104, S => n1032, Z => n2896);
   U879 : MUX2_X1 port map( A => n3813, B => n1105, S => n1032, Z => n2895);
   U880 : MUX2_X1 port map( A => n3812, B => n1106, S => n1032, Z => n2894);
   U881 : MUX2_X1 port map( A => n3811, B => n1107, S => n1032, Z => n2893);
   U882 : MUX2_X1 port map( A => n3810, B => n1108, S => n1032, Z => n2892);
   U883 : MUX2_X1 port map( A => n3809, B => n1109, S => n1032, Z => n2891);
   U884 : MUX2_X1 port map( A => n3808, B => n1110, S => n1032, Z => n2890);
   U885 : MUX2_X1 port map( A => n3807, B => n1111, S => n1032, Z => n2889);
   U886 : MUX2_X1 port map( A => n3806, B => n1112, S => n1032, Z => n2888);
   U887 : MUX2_X1 port map( A => n3805, B => n1113, S => n1032, Z => n2887);
   U888 : MUX2_X1 port map( A => n3804, B => n1114, S => n1032, Z => n2886);
   U889 : MUX2_X1 port map( A => n3803, B => n1115, S => n1032, Z => n2885);
   U890 : MUX2_X1 port map( A => n3802, B => n1116, S => n1032, Z => n2884);
   U891 : MUX2_X1 port map( A => n3801, B => n1117, S => n1032, Z => n2883);
   U892 : MUX2_X1 port map( A => n3800, B => n1118, S => n1032, Z => n2882);
   U893 : MUX2_X1 port map( A => n3799, B => n1119, S => n1032, Z => n2881);
   U894 : MUX2_X1 port map( A => n3798, B => n1120, S => n1032, Z => n2880);
   U895 : MUX2_X1 port map( A => n3797, B => n1121, S => n1032, Z => n2879);
   U896 : OAI21_X1 port map( B1 => n1135, B2 => n1150, A => RST, ZN => n1156);
   U897 : MUX2_X1 port map( A => n3796, B => n1089, S => n1034, Z => n2878);
   U898 : MUX2_X1 port map( A => n3795, B => n1091, S => n1034, Z => n2877);
   U899 : MUX2_X1 port map( A => n3794, B => n1092, S => n1034, Z => n2876);
   U900 : MUX2_X1 port map( A => n3793, B => n1093, S => n1034, Z => n2875);
   U901 : MUX2_X1 port map( A => n3792, B => n1094, S => n1034, Z => n2874);
   U902 : MUX2_X1 port map( A => n3791, B => n1095, S => n1034, Z => n2873);
   U903 : MUX2_X1 port map( A => n3790, B => n1096, S => n1034, Z => n2872);
   U904 : MUX2_X1 port map( A => n3789, B => n1097, S => n1034, Z => n2871);
   U905 : MUX2_X1 port map( A => n3788, B => n1098, S => n1034, Z => n2870);
   U906 : MUX2_X1 port map( A => n3787, B => n1099, S => n1034, Z => n2869);
   U907 : MUX2_X1 port map( A => n3786, B => n1100, S => n1034, Z => n2868);
   U908 : MUX2_X1 port map( A => n3785, B => n1101, S => n1034, Z => n2867);
   U909 : MUX2_X1 port map( A => n3784, B => n1102, S => n1034, Z => n2866);
   U910 : MUX2_X1 port map( A => n3783, B => n1103, S => n1034, Z => n2865);
   U911 : MUX2_X1 port map( A => n3782, B => n1104, S => n1034, Z => n2864);
   U912 : MUX2_X1 port map( A => n3781, B => n1105, S => n1034, Z => n2863);
   U913 : MUX2_X1 port map( A => n3780, B => n1106, S => n1034, Z => n2862);
   U914 : MUX2_X1 port map( A => n3779, B => n1107, S => n1034, Z => n2861);
   U915 : MUX2_X1 port map( A => n3778, B => n1108, S => n1034, Z => n2860);
   U916 : MUX2_X1 port map( A => n3777, B => n1109, S => n1034, Z => n2859);
   U917 : MUX2_X1 port map( A => n3776, B => n1110, S => n1034, Z => n2858);
   U918 : MUX2_X1 port map( A => n3775, B => n1111, S => n1034, Z => n2857);
   U919 : MUX2_X1 port map( A => n3774, B => n1112, S => n1034, Z => n2856);
   U920 : MUX2_X1 port map( A => n3773, B => n1113, S => n1034, Z => n2855);
   U921 : MUX2_X1 port map( A => n3772, B => n1114, S => n1034, Z => n2854);
   U922 : MUX2_X1 port map( A => n3771, B => n1115, S => n1034, Z => n2853);
   U923 : MUX2_X1 port map( A => n3770, B => n1116, S => n1034, Z => n2852);
   U924 : MUX2_X1 port map( A => n3769, B => n1117, S => n1034, Z => n2851);
   U925 : MUX2_X1 port map( A => n3768, B => n1118, S => n1034, Z => n2850);
   U926 : MUX2_X1 port map( A => n3767, B => n1119, S => n1034, Z => n2849);
   U927 : MUX2_X1 port map( A => n3766, B => n1120, S => n1034, Z => n2848);
   U928 : MUX2_X1 port map( A => n3765, B => n1121, S => n1034, Z => n2847);
   U929 : OAI21_X1 port map( B1 => n1137, B2 => n1150, A => RST, ZN => n1157);
   U930 : NAND3_X1 port map( A1 => WR, A2 => n1138, A3 => ADD_WR(4), ZN => 
                           n1150);
   U931 : INV_X1 port map( A => ADD_WR(3), ZN => n1138);
   U932 : MUX2_X1 port map( A => n3764, B => n1089, S => n1036, Z => n2846);
   U933 : MUX2_X1 port map( A => n3763, B => n1091, S => n1036, Z => n2845);
   U934 : MUX2_X1 port map( A => n3762, B => n1092, S => n1036, Z => n2844);
   U935 : MUX2_X1 port map( A => n3761, B => n1093, S => n1036, Z => n2843);
   U936 : MUX2_X1 port map( A => n3760, B => n1094, S => n1036, Z => n2842);
   U937 : MUX2_X1 port map( A => n3759, B => n1095, S => n1036, Z => n2841);
   U938 : MUX2_X1 port map( A => n3758, B => n1096, S => n1036, Z => n2840);
   U939 : MUX2_X1 port map( A => n3757, B => n1097, S => n1036, Z => n2839);
   U940 : MUX2_X1 port map( A => n3756, B => n1098, S => n1036, Z => n2838);
   U941 : MUX2_X1 port map( A => n3755, B => n1099, S => n1036, Z => n2837);
   U942 : MUX2_X1 port map( A => n3754, B => n1100, S => n1036, Z => n2836);
   U943 : MUX2_X1 port map( A => n3753, B => n1101, S => n1036, Z => n2835);
   U944 : MUX2_X1 port map( A => n3752, B => n1102, S => n1036, Z => n2834);
   U945 : MUX2_X1 port map( A => n3751, B => n1103, S => n1036, Z => n2833);
   U946 : MUX2_X1 port map( A => n3750, B => n1104, S => n1036, Z => n2832);
   U947 : MUX2_X1 port map( A => n3749, B => n1105, S => n1036, Z => n2831);
   U948 : MUX2_X1 port map( A => n3748, B => n1106, S => n1036, Z => n2830);
   U949 : MUX2_X1 port map( A => n3747, B => n1107, S => n1036, Z => n2829);
   U950 : MUX2_X1 port map( A => n3746, B => n1108, S => n1036, Z => n2828);
   U951 : MUX2_X1 port map( A => n3745, B => n1109, S => n1036, Z => n2827);
   U952 : MUX2_X1 port map( A => n3744, B => n1110, S => n1036, Z => n2826);
   U953 : MUX2_X1 port map( A => n3743, B => n1111, S => n1036, Z => n2825);
   U954 : MUX2_X1 port map( A => n3742, B => n1112, S => n1036, Z => n2824);
   U955 : MUX2_X1 port map( A => n3741, B => n1113, S => n1036, Z => n2823);
   U956 : MUX2_X1 port map( A => n3740, B => n1114, S => n1036, Z => n2822);
   U957 : MUX2_X1 port map( A => n3739, B => n1115, S => n1036, Z => n2821);
   U958 : MUX2_X1 port map( A => n3738, B => n1116, S => n1036, Z => n2820);
   U959 : MUX2_X1 port map( A => n3737, B => n1117, S => n1036, Z => n2819);
   U960 : MUX2_X1 port map( A => n3736, B => n1118, S => n1036, Z => n2818);
   U961 : MUX2_X1 port map( A => n3735, B => n1119, S => n1036, Z => n2817);
   U962 : MUX2_X1 port map( A => n3734, B => n1120, S => n1036, Z => n2816);
   U963 : MUX2_X1 port map( A => n3733, B => n1121, S => n1036, Z => n2815);
   U964 : OAI21_X1 port map( B1 => n1123, B2 => n1159, A => RST, ZN => n1158);
   U965 : NAND3_X1 port map( A1 => n1160, A2 => n1161, A3 => n1162, ZN => n1123
                           );
   U966 : MUX2_X1 port map( A => n3732, B => n1089, S => n1038, Z => n2814);
   U967 : MUX2_X1 port map( A => n3731, B => n1091, S => n1038, Z => n2813);
   U968 : MUX2_X1 port map( A => n3730, B => n1092, S => n1038, Z => n2812);
   U969 : MUX2_X1 port map( A => n3729, B => n1093, S => n1038, Z => n2811);
   U970 : MUX2_X1 port map( A => n3728, B => n1094, S => n1038, Z => n2810);
   U971 : MUX2_X1 port map( A => n3727, B => n1095, S => n1038, Z => n2809);
   U972 : MUX2_X1 port map( A => n3726, B => n1096, S => n1038, Z => n2808);
   U973 : MUX2_X1 port map( A => n3725, B => n1097, S => n1038, Z => n2807);
   U974 : MUX2_X1 port map( A => n3724, B => n1098, S => n1038, Z => n2806);
   U975 : MUX2_X1 port map( A => n3723, B => n1099, S => n1038, Z => n2805);
   U976 : MUX2_X1 port map( A => n3722, B => n1100, S => n1038, Z => n2804);
   U977 : MUX2_X1 port map( A => n3721, B => n1101, S => n1038, Z => n2803);
   U978 : MUX2_X1 port map( A => n3720, B => n1102, S => n1038, Z => n2802);
   U979 : MUX2_X1 port map( A => n3719, B => n1103, S => n1038, Z => n2801);
   U980 : MUX2_X1 port map( A => n3718, B => n1104, S => n1038, Z => n2800);
   U981 : MUX2_X1 port map( A => n3717, B => n1105, S => n1038, Z => n2799);
   U982 : MUX2_X1 port map( A => n3716, B => n1106, S => n1038, Z => n2798);
   U983 : MUX2_X1 port map( A => n3715, B => n1107, S => n1038, Z => n2797);
   U984 : MUX2_X1 port map( A => n3714, B => n1108, S => n1038, Z => n2796);
   U985 : MUX2_X1 port map( A => n3713, B => n1109, S => n1038, Z => n2795);
   U986 : MUX2_X1 port map( A => n3712, B => n1110, S => n1038, Z => n2794);
   U987 : MUX2_X1 port map( A => n3711, B => n1111, S => n1038, Z => n2793);
   U988 : MUX2_X1 port map( A => n3710, B => n1112, S => n1038, Z => n2792);
   U989 : MUX2_X1 port map( A => n3709, B => n1113, S => n1038, Z => n2791);
   U990 : MUX2_X1 port map( A => n3708, B => n1114, S => n1038, Z => n2790);
   U991 : MUX2_X1 port map( A => n3707, B => n1115, S => n1038, Z => n2789);
   U992 : MUX2_X1 port map( A => n3706, B => n1116, S => n1038, Z => n2788);
   U993 : MUX2_X1 port map( A => n3705, B => n1117, S => n1038, Z => n2787);
   U994 : MUX2_X1 port map( A => n3704, B => n1118, S => n1038, Z => n2786);
   U995 : MUX2_X1 port map( A => n3703, B => n1119, S => n1038, Z => n2785);
   U996 : MUX2_X1 port map( A => n3702, B => n1120, S => n1038, Z => n2784);
   U997 : MUX2_X1 port map( A => n3701, B => n1121, S => n1038, Z => n2783);
   U998 : OAI21_X1 port map( B1 => n1125, B2 => n1159, A => RST, ZN => n1163);
   U999 : NAND3_X1 port map( A1 => n1160, A2 => n1161, A3 => ADD_WR(0), ZN => 
                           n1125);
   U1000 : MUX2_X1 port map( A => n897, B => n1089, S => n1040, Z => n2782);
   U1001 : MUX2_X1 port map( A => n898, B => n1091, S => n1040, Z => n2781);
   U1002 : MUX2_X1 port map( A => n899, B => n1092, S => n1040, Z => n2780);
   U1003 : MUX2_X1 port map( A => n900, B => n1093, S => n1040, Z => n2779);
   U1004 : MUX2_X1 port map( A => n901, B => n1094, S => n1040, Z => n2778);
   U1005 : MUX2_X1 port map( A => n902, B => n1095, S => n1040, Z => n2777);
   U1006 : MUX2_X1 port map( A => n903, B => n1096, S => n1040, Z => n2776);
   U1007 : MUX2_X1 port map( A => n904, B => n1097, S => n1040, Z => n2775);
   U1008 : MUX2_X1 port map( A => n905, B => n1098, S => n1040, Z => n2774);
   U1009 : MUX2_X1 port map( A => n906, B => n1099, S => n1040, Z => n2773);
   U1010 : MUX2_X1 port map( A => n907, B => n1100, S => n1040, Z => n2772);
   U1011 : MUX2_X1 port map( A => n908, B => n1101, S => n1040, Z => n2771);
   U1012 : MUX2_X1 port map( A => n909, B => n1102, S => n1040, Z => n2770);
   U1013 : MUX2_X1 port map( A => n910, B => n1103, S => n1040, Z => n2769);
   U1014 : MUX2_X1 port map( A => n911, B => n1104, S => n1040, Z => n2768);
   U1015 : MUX2_X1 port map( A => n912, B => n1105, S => n1040, Z => n2767);
   U1016 : MUX2_X1 port map( A => n913, B => n1106, S => n1040, Z => n2766);
   U1017 : MUX2_X1 port map( A => n914, B => n1107, S => n1040, Z => n2765);
   U1018 : MUX2_X1 port map( A => n915, B => n1108, S => n1040, Z => n2764);
   U1019 : MUX2_X1 port map( A => n916, B => n1109, S => n1040, Z => n2763);
   U1020 : MUX2_X1 port map( A => n917, B => n1110, S => n1040, Z => n2762);
   U1021 : MUX2_X1 port map( A => n918, B => n1111, S => n1040, Z => n2761);
   U1022 : MUX2_X1 port map( A => n919, B => n1112, S => n1040, Z => n2760);
   U1023 : MUX2_X1 port map( A => n920, B => n1113, S => n1040, Z => n2759);
   U1024 : MUX2_X1 port map( A => n921, B => n1114, S => n1040, Z => n2758);
   U1025 : MUX2_X1 port map( A => n922, B => n1115, S => n1040, Z => n2757);
   U1026 : MUX2_X1 port map( A => n923, B => n1116, S => n1040, Z => n2756);
   U1027 : MUX2_X1 port map( A => n924, B => n1117, S => n1040, Z => n2755);
   U1028 : MUX2_X1 port map( A => n925, B => n1118, S => n1040, Z => n2754);
   U1029 : MUX2_X1 port map( A => n926, B => n1119, S => n1040, Z => n2753);
   U1030 : MUX2_X1 port map( A => n927, B => n1120, S => n1040, Z => n2752);
   U1031 : MUX2_X1 port map( A => n928, B => n1121, S => n1040, Z => n2751);
   U1032 : OAI21_X1 port map( B1 => n1127, B2 => n1159, A => RST, ZN => n1164);
   U1033 : NAND3_X1 port map( A1 => n1162, A2 => n1161, A3 => ADD_WR(1), ZN => 
                           n1127);
   U1034 : MUX2_X1 port map( A => n577, B => n1089, S => n1042, Z => n2750);
   U1035 : MUX2_X1 port map( A => n578, B => n1091, S => n1042, Z => n2749);
   U1036 : MUX2_X1 port map( A => n579, B => n1092, S => n1042, Z => n2748);
   U1037 : MUX2_X1 port map( A => n580, B => n1093, S => n1042, Z => n2747);
   U1038 : MUX2_X1 port map( A => n581, B => n1094, S => n1042, Z => n2746);
   U1039 : MUX2_X1 port map( A => n582, B => n1095, S => n1042, Z => n2745);
   U1040 : MUX2_X1 port map( A => n583, B => n1096, S => n1042, Z => n2744);
   U1041 : MUX2_X1 port map( A => n584, B => n1097, S => n1042, Z => n2743);
   U1042 : MUX2_X1 port map( A => n585, B => n1098, S => n1042, Z => n2742);
   U1043 : MUX2_X1 port map( A => n586, B => n1099, S => n1042, Z => n2741);
   U1044 : MUX2_X1 port map( A => n587, B => n1100, S => n1042, Z => n2740);
   U1045 : MUX2_X1 port map( A => n588, B => n1101, S => n1042, Z => n2739);
   U1046 : MUX2_X1 port map( A => n589, B => n1102, S => n1042, Z => n2738);
   U1047 : MUX2_X1 port map( A => n590, B => n1103, S => n1042, Z => n2737);
   U1048 : MUX2_X1 port map( A => n591, B => n1104, S => n1042, Z => n2736);
   U1049 : MUX2_X1 port map( A => n592, B => n1105, S => n1042, Z => n2735);
   U1050 : MUX2_X1 port map( A => n593, B => n1106, S => n1042, Z => n2734);
   U1051 : MUX2_X1 port map( A => n594, B => n1107, S => n1042, Z => n2733);
   U1052 : MUX2_X1 port map( A => n595, B => n1108, S => n1042, Z => n2732);
   U1053 : MUX2_X1 port map( A => n596, B => n1109, S => n1042, Z => n2731);
   U1054 : MUX2_X1 port map( A => n597, B => n1110, S => n1042, Z => n2730);
   U1055 : MUX2_X1 port map( A => n598, B => n1111, S => n1042, Z => n2729);
   U1056 : MUX2_X1 port map( A => n599, B => n1112, S => n1042, Z => n2728);
   U1057 : MUX2_X1 port map( A => n600, B => n1113, S => n1042, Z => n2727);
   U1058 : MUX2_X1 port map( A => n601, B => n1114, S => n1042, Z => n2726);
   U1059 : MUX2_X1 port map( A => n602, B => n1115, S => n1042, Z => n2725);
   U1060 : MUX2_X1 port map( A => n603, B => n1116, S => n1042, Z => n2724);
   U1061 : MUX2_X1 port map( A => n604, B => n1117, S => n1042, Z => n2723);
   U1062 : MUX2_X1 port map( A => n605, B => n1118, S => n1042, Z => n2722);
   U1063 : MUX2_X1 port map( A => n606, B => n1119, S => n1042, Z => n2721);
   U1064 : MUX2_X1 port map( A => n607, B => n1120, S => n1042, Z => n2720);
   U1065 : MUX2_X1 port map( A => n608, B => n1121, S => n1042, Z => n2719);
   U1066 : OAI21_X1 port map( B1 => n1129, B2 => n1159, A => RST, ZN => n1165);
   U1067 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1161, A3 => ADD_WR(1), ZN
                           => n1129);
   U1068 : INV_X1 port map( A => ADD_WR(2), ZN => n1161);
   U1069 : MUX2_X1 port map( A => n3700, B => n1089, S => n1044, Z => n2718);
   U1070 : MUX2_X1 port map( A => n3699, B => n1091, S => n1044, Z => n2717);
   U1071 : MUX2_X1 port map( A => n3698, B => n1092, S => n1044, Z => n2716);
   U1072 : MUX2_X1 port map( A => n3697, B => n1093, S => n1044, Z => n2715);
   U1073 : MUX2_X1 port map( A => n3696, B => n1094, S => n1044, Z => n2714);
   U1074 : MUX2_X1 port map( A => n3695, B => n1095, S => n1044, Z => n2713);
   U1075 : MUX2_X1 port map( A => n3694, B => n1096, S => n1044, Z => n2712);
   U1076 : MUX2_X1 port map( A => n3693, B => n1097, S => n1044, Z => n2711);
   U1077 : MUX2_X1 port map( A => n3692, B => n1098, S => n1044, Z => n2710);
   U1078 : MUX2_X1 port map( A => n3691, B => n1099, S => n1044, Z => n2709);
   U1079 : MUX2_X1 port map( A => n3690, B => n1100, S => n1044, Z => n2708);
   U1080 : MUX2_X1 port map( A => n3689, B => n1101, S => n1044, Z => n2707);
   U1081 : MUX2_X1 port map( A => n3688, B => n1102, S => n1044, Z => n2706);
   U1082 : MUX2_X1 port map( A => n3687, B => n1103, S => n1044, Z => n2705);
   U1083 : MUX2_X1 port map( A => n3686, B => n1104, S => n1044, Z => n2704);
   U1084 : MUX2_X1 port map( A => n3685, B => n1105, S => n1044, Z => n2703);
   U1085 : MUX2_X1 port map( A => n3684, B => n1106, S => n1044, Z => n2702);
   U1086 : MUX2_X1 port map( A => n3683, B => n1107, S => n1044, Z => n2701);
   U1087 : MUX2_X1 port map( A => n3682, B => n1108, S => n1044, Z => n2700);
   U1088 : MUX2_X1 port map( A => n3681, B => n1109, S => n1044, Z => n2699);
   U1089 : MUX2_X1 port map( A => n3680, B => n1110, S => n1044, Z => n2698);
   U1090 : MUX2_X1 port map( A => n3679, B => n1111, S => n1044, Z => n2697);
   U1091 : MUX2_X1 port map( A => n3678, B => n1112, S => n1044, Z => n2696);
   U1092 : MUX2_X1 port map( A => n3677, B => n1113, S => n1044, Z => n2695);
   U1093 : MUX2_X1 port map( A => n3676, B => n1114, S => n1044, Z => n2694);
   U1094 : MUX2_X1 port map( A => n3675, B => n1115, S => n1044, Z => n2693);
   U1095 : MUX2_X1 port map( A => n3674, B => n1116, S => n1044, Z => n2692);
   U1096 : MUX2_X1 port map( A => n3673, B => n1117, S => n1044, Z => n2691);
   U1097 : MUX2_X1 port map( A => n3672, B => n1118, S => n1044, Z => n2690);
   U1098 : MUX2_X1 port map( A => n3671, B => n1119, S => n1044, Z => n2689);
   U1099 : MUX2_X1 port map( A => n3670, B => n1120, S => n1044, Z => n2688);
   U1100 : MUX2_X1 port map( A => n3669, B => n1121, S => n1044, Z => n2687);
   U1101 : OAI21_X1 port map( B1 => n1131, B2 => n1159, A => RST, ZN => n1166);
   U1102 : NAND3_X1 port map( A1 => n1162, A2 => n1160, A3 => ADD_WR(2), ZN => 
                           n1131);
   U1103 : MUX2_X1 port map( A => n3668, B => n1089, S => n1046, Z => n2686);
   U1104 : MUX2_X1 port map( A => n3667, B => n1091, S => n1046, Z => n2685);
   U1105 : MUX2_X1 port map( A => n3666, B => n1092, S => n1046, Z => n2684);
   U1106 : MUX2_X1 port map( A => n3665, B => n1093, S => n1046, Z => n2683);
   U1107 : MUX2_X1 port map( A => n3664, B => n1094, S => n1046, Z => n2682);
   U1108 : MUX2_X1 port map( A => n3663, B => n1095, S => n1046, Z => n2681);
   U1109 : MUX2_X1 port map( A => n3662, B => n1096, S => n1046, Z => n2680);
   U1110 : MUX2_X1 port map( A => n3661, B => n1097, S => n1046, Z => n2679);
   U1111 : MUX2_X1 port map( A => n3660, B => n1098, S => n1046, Z => n2678);
   U1112 : MUX2_X1 port map( A => n3659, B => n1099, S => n1046, Z => n2677);
   U1113 : MUX2_X1 port map( A => n3658, B => n1100, S => n1046, Z => n2676);
   U1114 : MUX2_X1 port map( A => n3657, B => n1101, S => n1046, Z => n2675);
   U1115 : MUX2_X1 port map( A => n3656, B => n1102, S => n1046, Z => n2674);
   U1116 : MUX2_X1 port map( A => n3655, B => n1103, S => n1046, Z => n2673);
   U1117 : MUX2_X1 port map( A => n3654, B => n1104, S => n1046, Z => n2672);
   U1118 : MUX2_X1 port map( A => n3653, B => n1105, S => n1046, Z => n2671);
   U1119 : MUX2_X1 port map( A => n3652, B => n1106, S => n1046, Z => n2670);
   U1120 : MUX2_X1 port map( A => n3651, B => n1107, S => n1046, Z => n2669);
   U1121 : MUX2_X1 port map( A => n3650, B => n1108, S => n1046, Z => n2668);
   U1122 : MUX2_X1 port map( A => n3649, B => n1109, S => n1046, Z => n2667);
   U1123 : MUX2_X1 port map( A => n3648, B => n1110, S => n1046, Z => n2666);
   U1124 : MUX2_X1 port map( A => n3647, B => n1111, S => n1046, Z => n2665);
   U1125 : MUX2_X1 port map( A => n3646, B => n1112, S => n1046, Z => n2664);
   U1126 : MUX2_X1 port map( A => n3645, B => n1113, S => n1046, Z => n2663);
   U1127 : MUX2_X1 port map( A => n3644, B => n1114, S => n1046, Z => n2662);
   U1128 : MUX2_X1 port map( A => n3643, B => n1115, S => n1046, Z => n2661);
   U1129 : MUX2_X1 port map( A => n3642, B => n1116, S => n1046, Z => n2660);
   U1130 : MUX2_X1 port map( A => n3641, B => n1117, S => n1046, Z => n2659);
   U1131 : MUX2_X1 port map( A => n3640, B => n1118, S => n1046, Z => n2658);
   U1132 : MUX2_X1 port map( A => n3639, B => n1119, S => n1046, Z => n2657);
   U1133 : MUX2_X1 port map( A => n3638, B => n1120, S => n1046, Z => n2656);
   U1134 : MUX2_X1 port map( A => n3637, B => n1121, S => n1046, Z => n2655);
   U1135 : OAI21_X1 port map( B1 => n1133, B2 => n1159, A => RST, ZN => n1167);
   U1136 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1160, A3 => ADD_WR(2), ZN
                           => n1133);
   U1137 : INV_X1 port map( A => ADD_WR(1), ZN => n1160);
   U1138 : MUX2_X1 port map( A => n929, B => n1089, S => n1048, Z => n2654);
   U1139 : MUX2_X1 port map( A => n930, B => n1091, S => n1048, Z => n2653);
   U1140 : MUX2_X1 port map( A => n931, B => n1092, S => n1048, Z => n2652);
   U1141 : MUX2_X1 port map( A => n932, B => n1093, S => n1048, Z => n2651);
   U1142 : MUX2_X1 port map( A => n933, B => n1094, S => n1048, Z => n2650);
   U1143 : MUX2_X1 port map( A => n934, B => n1095, S => n1048, Z => n2649);
   U1144 : MUX2_X1 port map( A => n935, B => n1096, S => n1048, Z => n2648);
   U1145 : MUX2_X1 port map( A => n936, B => n1097, S => n1048, Z => n2647);
   U1146 : MUX2_X1 port map( A => n937, B => n1098, S => n1048, Z => n2646);
   U1147 : MUX2_X1 port map( A => n938, B => n1099, S => n1048, Z => n2645);
   U1148 : MUX2_X1 port map( A => n939, B => n1100, S => n1048, Z => n2644);
   U1149 : MUX2_X1 port map( A => n940, B => n1101, S => n1048, Z => n2643);
   U1150 : MUX2_X1 port map( A => n941, B => n1102, S => n1048, Z => n2642);
   U1151 : MUX2_X1 port map( A => n942, B => n1103, S => n1048, Z => n2641);
   U1152 : MUX2_X1 port map( A => n943, B => n1104, S => n1048, Z => n2640);
   U1153 : MUX2_X1 port map( A => n944, B => n1105, S => n1048, Z => n2639);
   U1154 : MUX2_X1 port map( A => n945, B => n1106, S => n1048, Z => n2638);
   U1155 : MUX2_X1 port map( A => n946, B => n1107, S => n1048, Z => n2637);
   U1156 : MUX2_X1 port map( A => n947, B => n1108, S => n1048, Z => n2636);
   U1157 : MUX2_X1 port map( A => n948, B => n1109, S => n1048, Z => n2635);
   U1158 : MUX2_X1 port map( A => n949, B => n1110, S => n1048, Z => n2634);
   U1159 : MUX2_X1 port map( A => n950, B => n1111, S => n1048, Z => n2633);
   U1160 : MUX2_X1 port map( A => n951, B => n1112, S => n1048, Z => n2632);
   U1161 : MUX2_X1 port map( A => n952, B => n1113, S => n1048, Z => n2631);
   U1162 : MUX2_X1 port map( A => n953, B => n1114, S => n1048, Z => n2630);
   U1163 : MUX2_X1 port map( A => n954, B => n1115, S => n1048, Z => n2629);
   U1164 : MUX2_X1 port map( A => n955, B => n1116, S => n1048, Z => n2628);
   U1165 : MUX2_X1 port map( A => n956, B => n1117, S => n1048, Z => n2627);
   U1166 : MUX2_X1 port map( A => n957, B => n1118, S => n1048, Z => n2626);
   U1167 : MUX2_X1 port map( A => n958, B => n1119, S => n1048, Z => n2625);
   U1168 : MUX2_X1 port map( A => n959, B => n1120, S => n1048, Z => n2624);
   U1169 : MUX2_X1 port map( A => n960, B => n1121, S => n1048, Z => n2623);
   U1170 : OAI21_X1 port map( B1 => n1135, B2 => n1159, A => RST, ZN => n1168);
   U1171 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n1162, A3 => ADD_WR(2), ZN
                           => n1135);
   U1172 : INV_X1 port map( A => ADD_WR(0), ZN => n1162);
   U1173 : MUX2_X1 port map( A => n609, B => n1089, S => n1050, Z => n2622);
   U1174 : AND2_X1 port map( A1 => RST, A2 => DATAIN(31), ZN => n1089);
   U1175 : MUX2_X1 port map( A => n610, B => n1091, S => n1050, Z => n2621);
   U1176 : AND2_X1 port map( A1 => DATAIN(30), A2 => RST, ZN => n1091);
   U1177 : MUX2_X1 port map( A => n611, B => n1092, S => n1050, Z => n2620);
   U1178 : AND2_X1 port map( A1 => DATAIN(29), A2 => RST, ZN => n1092);
   U1179 : MUX2_X1 port map( A => n612, B => n1093, S => n1050, Z => n2619);
   U1180 : AND2_X1 port map( A1 => DATAIN(28), A2 => RST, ZN => n1093);
   U1181 : MUX2_X1 port map( A => n613, B => n1094, S => n1050, Z => n2618);
   U1182 : AND2_X1 port map( A1 => DATAIN(27), A2 => RST, ZN => n1094);
   U1183 : MUX2_X1 port map( A => n614, B => n1095, S => n1050, Z => n2617);
   U1184 : AND2_X1 port map( A1 => DATAIN(26), A2 => RST, ZN => n1095);
   U1185 : MUX2_X1 port map( A => n615, B => n1096, S => n1050, Z => n2616);
   U1186 : AND2_X1 port map( A1 => DATAIN(25), A2 => RST, ZN => n1096);
   U1187 : MUX2_X1 port map( A => n616, B => n1097, S => n1050, Z => n2615);
   U1188 : AND2_X1 port map( A1 => DATAIN(24), A2 => RST, ZN => n1097);
   U1189 : MUX2_X1 port map( A => n617, B => n1098, S => n1050, Z => n2614);
   U1190 : AND2_X1 port map( A1 => DATAIN(23), A2 => RST, ZN => n1098);
   U1191 : MUX2_X1 port map( A => n618, B => n1099, S => n1050, Z => n2613);
   U1192 : AND2_X1 port map( A1 => DATAIN(22), A2 => RST, ZN => n1099);
   U1193 : MUX2_X1 port map( A => n619, B => n1100, S => n1050, Z => n2612);
   U1194 : AND2_X1 port map( A1 => DATAIN(21), A2 => RST, ZN => n1100);
   U1195 : MUX2_X1 port map( A => n620, B => n1101, S => n1050, Z => n2611);
   U1196 : AND2_X1 port map( A1 => DATAIN(20), A2 => RST, ZN => n1101);
   U1197 : MUX2_X1 port map( A => n621, B => n1102, S => n1050, Z => n2610);
   U1198 : AND2_X1 port map( A1 => DATAIN(19), A2 => RST, ZN => n1102);
   U1199 : MUX2_X1 port map( A => n622, B => n1103, S => n1050, Z => n2609);
   U1200 : AND2_X1 port map( A1 => DATAIN(18), A2 => RST, ZN => n1103);
   U1201 : MUX2_X1 port map( A => n623, B => n1104, S => n1050, Z => n2608);
   U1202 : AND2_X1 port map( A1 => DATAIN(17), A2 => RST, ZN => n1104);
   U1203 : MUX2_X1 port map( A => n624, B => n1105, S => n1050, Z => n2607);
   U1204 : AND2_X1 port map( A1 => DATAIN(16), A2 => RST, ZN => n1105);
   U1205 : MUX2_X1 port map( A => n625, B => n1106, S => n1050, Z => n2606);
   U1206 : AND2_X1 port map( A1 => DATAIN(15), A2 => RST, ZN => n1106);
   U1207 : MUX2_X1 port map( A => n626, B => n1107, S => n1050, Z => n2605);
   U1208 : AND2_X1 port map( A1 => DATAIN(14), A2 => RST, ZN => n1107);
   U1209 : MUX2_X1 port map( A => n627, B => n1108, S => n1050, Z => n2604);
   U1210 : AND2_X1 port map( A1 => DATAIN(13), A2 => RST, ZN => n1108);
   U1211 : MUX2_X1 port map( A => n628, B => n1109, S => n1050, Z => n2603);
   U1212 : AND2_X1 port map( A1 => DATAIN(12), A2 => RST, ZN => n1109);
   U1213 : MUX2_X1 port map( A => n629, B => n1110, S => n1050, Z => n2602);
   U1214 : AND2_X1 port map( A1 => DATAIN(11), A2 => RST, ZN => n1110);
   U1215 : MUX2_X1 port map( A => n630, B => n1111, S => n1050, Z => n2601);
   U1216 : AND2_X1 port map( A1 => DATAIN(10), A2 => RST, ZN => n1111);
   U1217 : MUX2_X1 port map( A => n631, B => n1112, S => n1050, Z => n2600);
   U1218 : AND2_X1 port map( A1 => DATAIN(9), A2 => RST, ZN => n1112);
   U1219 : MUX2_X1 port map( A => n632, B => n1113, S => n1050, Z => n2599);
   U1220 : AND2_X1 port map( A1 => DATAIN(8), A2 => RST, ZN => n1113);
   U1221 : MUX2_X1 port map( A => n633, B => n1114, S => n1050, Z => n2598);
   U1222 : AND2_X1 port map( A1 => DATAIN(7), A2 => RST, ZN => n1114);
   U1223 : MUX2_X1 port map( A => n634, B => n1115, S => n1050, Z => n2597);
   U1224 : AND2_X1 port map( A1 => DATAIN(6), A2 => RST, ZN => n1115);
   U1225 : MUX2_X1 port map( A => n635, B => n1116, S => n1050, Z => n2596);
   U1226 : AND2_X1 port map( A1 => DATAIN(5), A2 => RST, ZN => n1116);
   U1227 : MUX2_X1 port map( A => n636, B => n1117, S => n1050, Z => n2595);
   U1228 : AND2_X1 port map( A1 => DATAIN(4), A2 => RST, ZN => n1117);
   U1229 : MUX2_X1 port map( A => n637, B => n1118, S => n1050, Z => n2594);
   U1230 : AND2_X1 port map( A1 => DATAIN(3), A2 => RST, ZN => n1118);
   U1231 : MUX2_X1 port map( A => n638, B => n1119, S => n1050, Z => n2593);
   U1232 : AND2_X1 port map( A1 => DATAIN(2), A2 => RST, ZN => n1119);
   U1233 : MUX2_X1 port map( A => n639, B => n1120, S => n1050, Z => n2592);
   U1234 : AND2_X1 port map( A1 => DATAIN(1), A2 => RST, ZN => n1120);
   U1235 : MUX2_X1 port map( A => n640, B => n1121, S => n1050, Z => n2591);
   U1236 : OAI21_X1 port map( B1 => n1137, B2 => n1159, A => RST, ZN => n1169);
   U1237 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => WR, A3 => ADD_WR(4), ZN =>
                           n1159);
   U1238 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n1137);
   U1239 : AND2_X1 port map( A1 => DATAIN(0), A2 => RST, ZN => n1121);
   U1240 : OAI22_X1 port map( A1 => n3636, A2 => n1170, B1 => n1171, B2 => 
                           n1172, ZN => n2590);
   U1241 : NOR2_X1 port map( A1 => n1173, A2 => n1174, ZN => n1171);
   U1242 : NAND4_X1 port map( A1 => n1175, A2 => n1176, A3 => n1177, A4 => 
                           n1178, ZN => n1174);
   U1243 : AOI221_X1 port map( B1 => n1179, B2 => n3668, C1 => n1180, C2 => 
                           n3700, A => n1181, ZN => n1178);
   U1244 : OAI22_X1 port map( A1 => n993, A2 => n1182, B1 => n961, B2 => n1183,
                           ZN => n1181);
   U1245 : AOI221_X1 port map( B1 => n1184, B2 => n3732, C1 => n1185, C2 => 
                           n3764, A => n1186, ZN => n1177);
   U1246 : OAI22_X1 port map( A1 => n865, A2 => n1187, B1 => n833, B2 => n1188,
                           ZN => n1186);
   U1247 : AOI221_X1 port map( B1 => n1189, B2 => n3796, C1 => n1190, C2 => 
                           n3828, A => n1191, ZN => n1176);
   U1248 : OAI22_X1 port map( A1 => n673, A2 => n1192, B1 => n641, B2 => n1193,
                           ZN => n1191);
   U1249 : AOI221_X1 port map( B1 => n1194, B2 => n3860, C1 => n1195, C2 => 
                           n3892, A => n1196, ZN => n1175);
   U1250 : OAI22_X1 port map( A1 => n545, A2 => n1197, B1 => n513, B2 => n1198,
                           ZN => n1196);
   U1251 : NAND4_X1 port map( A1 => n1199, A2 => n1200, A3 => n1201, A4 => 
                           n1202, ZN => n1173);
   U1252 : AOI221_X1 port map( B1 => n1203, B2 => n3924, C1 => n1204, C2 => 
                           n3956, A => n1205, ZN => n1202);
   U1253 : OAI22_X1 port map( A1 => n417, A2 => n1206, B1 => n385, B2 => n1207,
                           ZN => n1205);
   U1254 : AOI221_X1 port map( B1 => n1208, B2 => n3988, C1 => n1209, C2 => 
                           n4020, A => n1210, ZN => n1201);
   U1255 : OAI22_X1 port map( A1 => n289, A2 => n1211, B1 => n257, B2 => n1212,
                           ZN => n1210);
   U1256 : AOI221_X1 port map( B1 => n1213, B2 => n129, C1 => n1214, C2 => n1, 
                           A => n1215, ZN => n1200);
   U1257 : OAI22_X1 port map( A1 => n65, A2 => n1216, B1 => n193, B2 => n1217, 
                           ZN => n1215);
   U1258 : AOI221_X1 port map( B1 => n1218, B2 => n130, C1 => n1219, C2 => n2, 
                           A => n1220, ZN => n1199);
   U1259 : OAI22_X1 port map( A1 => n66, A2 => n1221, B1 => n194, B2 => n1222, 
                           ZN => n1220);
   U1260 : OAI22_X1 port map( A1 => n3635, A2 => n1170, B1 => n1223, B2 => 
                           n1172, ZN => n2589);
   U1261 : NOR2_X1 port map( A1 => n1224, A2 => n1225, ZN => n1223);
   U1262 : NAND4_X1 port map( A1 => n1226, A2 => n1227, A3 => n1228, A4 => 
                           n1229, ZN => n1225);
   U1263 : AOI221_X1 port map( B1 => n1179, B2 => n3667, C1 => n1180, C2 => 
                           n3699, A => n1230, ZN => n1229);
   U1264 : OAI22_X1 port map( A1 => n994, A2 => n1182, B1 => n962, B2 => n1183,
                           ZN => n1230);
   U1265 : AOI221_X1 port map( B1 => n1184, B2 => n3731, C1 => n1185, C2 => 
                           n3763, A => n1231, ZN => n1228);
   U1266 : OAI22_X1 port map( A1 => n866, A2 => n1187, B1 => n834, B2 => n1188,
                           ZN => n1231);
   U1267 : AOI221_X1 port map( B1 => n1189, B2 => n3795, C1 => n1190, C2 => 
                           n3827, A => n1232, ZN => n1227);
   U1268 : OAI22_X1 port map( A1 => n674, A2 => n1192, B1 => n642, B2 => n1193,
                           ZN => n1232);
   U1269 : AOI221_X1 port map( B1 => n1194, B2 => n3859, C1 => n1195, C2 => 
                           n3891, A => n1233, ZN => n1226);
   U1270 : OAI22_X1 port map( A1 => n546, A2 => n1197, B1 => n514, B2 => n1198,
                           ZN => n1233);
   U1271 : NAND4_X1 port map( A1 => n1234, A2 => n1235, A3 => n1236, A4 => 
                           n1237, ZN => n1224);
   U1272 : AOI221_X1 port map( B1 => n1203, B2 => n3923, C1 => n1204, C2 => 
                           n3955, A => n1238, ZN => n1237);
   U1273 : OAI22_X1 port map( A1 => n418, A2 => n1206, B1 => n386, B2 => n1207,
                           ZN => n1238);
   U1274 : AOI221_X1 port map( B1 => n1208, B2 => n3987, C1 => n1209, C2 => 
                           n4019, A => n1239, ZN => n1236);
   U1275 : OAI22_X1 port map( A1 => n290, A2 => n1211, B1 => n258, B2 => n1212,
                           ZN => n1239);
   U1276 : AOI221_X1 port map( B1 => n1213, B2 => n131, C1 => n1214, C2 => n3, 
                           A => n1240, ZN => n1235);
   U1277 : OAI22_X1 port map( A1 => n67, A2 => n1216, B1 => n195, B2 => n1217, 
                           ZN => n1240);
   U1278 : AOI221_X1 port map( B1 => n1218, B2 => n132, C1 => n1219, C2 => n4, 
                           A => n1241, ZN => n1234);
   U1279 : OAI22_X1 port map( A1 => n68, A2 => n1221, B1 => n196, B2 => n1222, 
                           ZN => n1241);
   U1280 : OAI22_X1 port map( A1 => n3634, A2 => n1170, B1 => n1242, B2 => 
                           n1172, ZN => n2588);
   U1281 : NOR2_X1 port map( A1 => n1243, A2 => n1244, ZN => n1242);
   U1282 : NAND4_X1 port map( A1 => n1245, A2 => n1246, A3 => n1247, A4 => 
                           n1248, ZN => n1244);
   U1283 : AOI221_X1 port map( B1 => n1179, B2 => n3666, C1 => n1180, C2 => 
                           n3698, A => n1249, ZN => n1248);
   U1284 : OAI22_X1 port map( A1 => n995, A2 => n1182, B1 => n963, B2 => n1183,
                           ZN => n1249);
   U1285 : AOI221_X1 port map( B1 => n1184, B2 => n3730, C1 => n1185, C2 => 
                           n3762, A => n1250, ZN => n1247);
   U1286 : OAI22_X1 port map( A1 => n867, A2 => n1187, B1 => n835, B2 => n1188,
                           ZN => n1250);
   U1287 : AOI221_X1 port map( B1 => n1189, B2 => n3794, C1 => n1190, C2 => 
                           n3826, A => n1251, ZN => n1246);
   U1288 : OAI22_X1 port map( A1 => n675, A2 => n1192, B1 => n643, B2 => n1193,
                           ZN => n1251);
   U1289 : AOI221_X1 port map( B1 => n1194, B2 => n3858, C1 => n1195, C2 => 
                           n3890, A => n1252, ZN => n1245);
   U1290 : OAI22_X1 port map( A1 => n547, A2 => n1197, B1 => n515, B2 => n1198,
                           ZN => n1252);
   U1291 : NAND4_X1 port map( A1 => n1253, A2 => n1254, A3 => n1255, A4 => 
                           n1256, ZN => n1243);
   U1292 : AOI221_X1 port map( B1 => n1203, B2 => n3922, C1 => n1204, C2 => 
                           n3954, A => n1257, ZN => n1256);
   U1293 : OAI22_X1 port map( A1 => n419, A2 => n1206, B1 => n387, B2 => n1207,
                           ZN => n1257);
   U1294 : AOI221_X1 port map( B1 => n1208, B2 => n3986, C1 => n1209, C2 => 
                           n4018, A => n1258, ZN => n1255);
   U1295 : OAI22_X1 port map( A1 => n291, A2 => n1211, B1 => n259, B2 => n1212,
                           ZN => n1258);
   U1296 : AOI221_X1 port map( B1 => n1213, B2 => n133, C1 => n1214, C2 => n5, 
                           A => n1259, ZN => n1254);
   U1297 : OAI22_X1 port map( A1 => n69, A2 => n1216, B1 => n197, B2 => n1217, 
                           ZN => n1259);
   U1298 : AOI221_X1 port map( B1 => n1218, B2 => n134, C1 => n1219, C2 => n6, 
                           A => n1260, ZN => n1253);
   U1299 : OAI22_X1 port map( A1 => n70, A2 => n1221, B1 => n198, B2 => n1222, 
                           ZN => n1260);
   U1300 : OAI22_X1 port map( A1 => n3633, A2 => n1170, B1 => n1261, B2 => 
                           n1172, ZN => n2587);
   U1301 : NOR2_X1 port map( A1 => n1262, A2 => n1263, ZN => n1261);
   U1302 : NAND4_X1 port map( A1 => n1264, A2 => n1265, A3 => n1266, A4 => 
                           n1267, ZN => n1263);
   U1303 : AOI221_X1 port map( B1 => n1179, B2 => n3665, C1 => n1180, C2 => 
                           n3697, A => n1268, ZN => n1267);
   U1304 : OAI22_X1 port map( A1 => n996, A2 => n1182, B1 => n964, B2 => n1183,
                           ZN => n1268);
   U1305 : AOI221_X1 port map( B1 => n1184, B2 => n3729, C1 => n1185, C2 => 
                           n3761, A => n1269, ZN => n1266);
   U1306 : OAI22_X1 port map( A1 => n868, A2 => n1187, B1 => n836, B2 => n1188,
                           ZN => n1269);
   U1307 : AOI221_X1 port map( B1 => n1189, B2 => n3793, C1 => n1190, C2 => 
                           n3825, A => n1270, ZN => n1265);
   U1308 : OAI22_X1 port map( A1 => n676, A2 => n1192, B1 => n644, B2 => n1193,
                           ZN => n1270);
   U1309 : AOI221_X1 port map( B1 => n1194, B2 => n3857, C1 => n1195, C2 => 
                           n3889, A => n1271, ZN => n1264);
   U1310 : OAI22_X1 port map( A1 => n548, A2 => n1197, B1 => n516, B2 => n1198,
                           ZN => n1271);
   U1311 : NAND4_X1 port map( A1 => n1272, A2 => n1273, A3 => n1274, A4 => 
                           n1275, ZN => n1262);
   U1312 : AOI221_X1 port map( B1 => n1203, B2 => n3921, C1 => n1204, C2 => 
                           n3953, A => n1276, ZN => n1275);
   U1313 : OAI22_X1 port map( A1 => n420, A2 => n1206, B1 => n388, B2 => n1207,
                           ZN => n1276);
   U1314 : AOI221_X1 port map( B1 => n1208, B2 => n3985, C1 => n1209, C2 => 
                           n4017, A => n1277, ZN => n1274);
   U1315 : OAI22_X1 port map( A1 => n292, A2 => n1211, B1 => n260, B2 => n1212,
                           ZN => n1277);
   U1316 : AOI221_X1 port map( B1 => n1213, B2 => n135, C1 => n1214, C2 => n7, 
                           A => n1278, ZN => n1273);
   U1317 : OAI22_X1 port map( A1 => n71, A2 => n1216, B1 => n199, B2 => n1217, 
                           ZN => n1278);
   U1318 : AOI221_X1 port map( B1 => n1218, B2 => n136, C1 => n1219, C2 => n8, 
                           A => n1279, ZN => n1272);
   U1319 : OAI22_X1 port map( A1 => n72, A2 => n1221, B1 => n200, B2 => n1222, 
                           ZN => n1279);
   U1320 : OAI22_X1 port map( A1 => n3632, A2 => n1170, B1 => n1280, B2 => 
                           n1172, ZN => n2586);
   U1321 : NOR2_X1 port map( A1 => n1281, A2 => n1282, ZN => n1280);
   U1322 : NAND4_X1 port map( A1 => n1283, A2 => n1284, A3 => n1285, A4 => 
                           n1286, ZN => n1282);
   U1323 : AOI221_X1 port map( B1 => n1179, B2 => n3664, C1 => n1180, C2 => 
                           n3696, A => n1287, ZN => n1286);
   U1324 : OAI22_X1 port map( A1 => n997, A2 => n1182, B1 => n965, B2 => n1183,
                           ZN => n1287);
   U1325 : AOI221_X1 port map( B1 => n1184, B2 => n3728, C1 => n1185, C2 => 
                           n3760, A => n1288, ZN => n1285);
   U1326 : OAI22_X1 port map( A1 => n869, A2 => n1187, B1 => n837, B2 => n1188,
                           ZN => n1288);
   U1327 : AOI221_X1 port map( B1 => n1189, B2 => n3792, C1 => n1190, C2 => 
                           n3824, A => n1289, ZN => n1284);
   U1328 : OAI22_X1 port map( A1 => n677, A2 => n1192, B1 => n645, B2 => n1193,
                           ZN => n1289);
   U1329 : AOI221_X1 port map( B1 => n1194, B2 => n3856, C1 => n1195, C2 => 
                           n3888, A => n1290, ZN => n1283);
   U1330 : OAI22_X1 port map( A1 => n549, A2 => n1197, B1 => n517, B2 => n1198,
                           ZN => n1290);
   U1331 : NAND4_X1 port map( A1 => n1291, A2 => n1292, A3 => n1293, A4 => 
                           n1294, ZN => n1281);
   U1332 : AOI221_X1 port map( B1 => n1203, B2 => n3920, C1 => n1204, C2 => 
                           n3952, A => n1295, ZN => n1294);
   U1333 : OAI22_X1 port map( A1 => n421, A2 => n1206, B1 => n389, B2 => n1207,
                           ZN => n1295);
   U1334 : AOI221_X1 port map( B1 => n1208, B2 => n3984, C1 => n1209, C2 => 
                           n4016, A => n1296, ZN => n1293);
   U1335 : OAI22_X1 port map( A1 => n293, A2 => n1211, B1 => n261, B2 => n1212,
                           ZN => n1296);
   U1336 : AOI221_X1 port map( B1 => n1213, B2 => n137, C1 => n1214, C2 => n9, 
                           A => n1297, ZN => n1292);
   U1337 : OAI22_X1 port map( A1 => n73, A2 => n1216, B1 => n201, B2 => n1217, 
                           ZN => n1297);
   U1338 : AOI221_X1 port map( B1 => n1218, B2 => n138, C1 => n1219, C2 => n10,
                           A => n1298, ZN => n1291);
   U1339 : OAI22_X1 port map( A1 => n74, A2 => n1221, B1 => n202, B2 => n1222, 
                           ZN => n1298);
   U1340 : OAI22_X1 port map( A1 => n3631, A2 => n1170, B1 => n1299, B2 => 
                           n1172, ZN => n2585);
   U1341 : NOR2_X1 port map( A1 => n1300, A2 => n1301, ZN => n1299);
   U1342 : NAND4_X1 port map( A1 => n1302, A2 => n1303, A3 => n1304, A4 => 
                           n1305, ZN => n1301);
   U1343 : AOI221_X1 port map( B1 => n1179, B2 => n3663, C1 => n1180, C2 => 
                           n3695, A => n1306, ZN => n1305);
   U1344 : OAI22_X1 port map( A1 => n998, A2 => n1182, B1 => n966, B2 => n1183,
                           ZN => n1306);
   U1345 : AOI221_X1 port map( B1 => n1184, B2 => n3727, C1 => n1185, C2 => 
                           n3759, A => n1307, ZN => n1304);
   U1346 : OAI22_X1 port map( A1 => n870, A2 => n1187, B1 => n838, B2 => n1188,
                           ZN => n1307);
   U1347 : AOI221_X1 port map( B1 => n1189, B2 => n3791, C1 => n1190, C2 => 
                           n3823, A => n1308, ZN => n1303);
   U1348 : OAI22_X1 port map( A1 => n678, A2 => n1192, B1 => n646, B2 => n1193,
                           ZN => n1308);
   U1349 : AOI221_X1 port map( B1 => n1194, B2 => n3855, C1 => n1195, C2 => 
                           n3887, A => n1309, ZN => n1302);
   U1350 : OAI22_X1 port map( A1 => n550, A2 => n1197, B1 => n518, B2 => n1198,
                           ZN => n1309);
   U1351 : NAND4_X1 port map( A1 => n1310, A2 => n1311, A3 => n1312, A4 => 
                           n1313, ZN => n1300);
   U1352 : AOI221_X1 port map( B1 => n1203, B2 => n3919, C1 => n1204, C2 => 
                           n3951, A => n1314, ZN => n1313);
   U1353 : OAI22_X1 port map( A1 => n422, A2 => n1206, B1 => n390, B2 => n1207,
                           ZN => n1314);
   U1354 : AOI221_X1 port map( B1 => n1208, B2 => n3983, C1 => n1209, C2 => 
                           n4015, A => n1315, ZN => n1312);
   U1355 : OAI22_X1 port map( A1 => n294, A2 => n1211, B1 => n262, B2 => n1212,
                           ZN => n1315);
   U1356 : AOI221_X1 port map( B1 => n1213, B2 => n139, C1 => n1214, C2 => n11,
                           A => n1316, ZN => n1311);
   U1357 : OAI22_X1 port map( A1 => n75, A2 => n1216, B1 => n203, B2 => n1217, 
                           ZN => n1316);
   U1358 : AOI221_X1 port map( B1 => n1218, B2 => n140, C1 => n1219, C2 => n12,
                           A => n1317, ZN => n1310);
   U1359 : OAI22_X1 port map( A1 => n76, A2 => n1221, B1 => n204, B2 => n1222, 
                           ZN => n1317);
   U1360 : OAI22_X1 port map( A1 => n3630, A2 => n1170, B1 => n1318, B2 => 
                           n1172, ZN => n2584);
   U1361 : NOR2_X1 port map( A1 => n1319, A2 => n1320, ZN => n1318);
   U1362 : NAND4_X1 port map( A1 => n1321, A2 => n1322, A3 => n1323, A4 => 
                           n1324, ZN => n1320);
   U1363 : AOI221_X1 port map( B1 => n1179, B2 => n3662, C1 => n1180, C2 => 
                           n3694, A => n1325, ZN => n1324);
   U1364 : OAI22_X1 port map( A1 => n999, A2 => n1182, B1 => n967, B2 => n1183,
                           ZN => n1325);
   U1365 : AOI221_X1 port map( B1 => n1184, B2 => n3726, C1 => n1185, C2 => 
                           n3758, A => n1326, ZN => n1323);
   U1366 : OAI22_X1 port map( A1 => n871, A2 => n1187, B1 => n839, B2 => n1188,
                           ZN => n1326);
   U1367 : AOI221_X1 port map( B1 => n1189, B2 => n3790, C1 => n1190, C2 => 
                           n3822, A => n1327, ZN => n1322);
   U1368 : OAI22_X1 port map( A1 => n679, A2 => n1192, B1 => n647, B2 => n1193,
                           ZN => n1327);
   U1369 : AOI221_X1 port map( B1 => n1194, B2 => n3854, C1 => n1195, C2 => 
                           n3886, A => n1328, ZN => n1321);
   U1370 : OAI22_X1 port map( A1 => n551, A2 => n1197, B1 => n519, B2 => n1198,
                           ZN => n1328);
   U1371 : NAND4_X1 port map( A1 => n1329, A2 => n1330, A3 => n1331, A4 => 
                           n1332, ZN => n1319);
   U1372 : AOI221_X1 port map( B1 => n1203, B2 => n3918, C1 => n1204, C2 => 
                           n3950, A => n1333, ZN => n1332);
   U1373 : OAI22_X1 port map( A1 => n423, A2 => n1206, B1 => n391, B2 => n1207,
                           ZN => n1333);
   U1374 : AOI221_X1 port map( B1 => n1208, B2 => n3982, C1 => n1209, C2 => 
                           n4014, A => n1334, ZN => n1331);
   U1375 : OAI22_X1 port map( A1 => n295, A2 => n1211, B1 => n263, B2 => n1212,
                           ZN => n1334);
   U1376 : AOI221_X1 port map( B1 => n1213, B2 => n141, C1 => n1214, C2 => n13,
                           A => n1335, ZN => n1330);
   U1377 : OAI22_X1 port map( A1 => n77, A2 => n1216, B1 => n205, B2 => n1217, 
                           ZN => n1335);
   U1378 : AOI221_X1 port map( B1 => n1218, B2 => n142, C1 => n1219, C2 => n14,
                           A => n1336, ZN => n1329);
   U1379 : OAI22_X1 port map( A1 => n78, A2 => n1221, B1 => n206, B2 => n1222, 
                           ZN => n1336);
   U1380 : OAI22_X1 port map( A1 => n3629, A2 => n1170, B1 => n1337, B2 => 
                           n1172, ZN => n2583);
   U1381 : NOR2_X1 port map( A1 => n1338, A2 => n1339, ZN => n1337);
   U1382 : NAND4_X1 port map( A1 => n1340, A2 => n1341, A3 => n1342, A4 => 
                           n1343, ZN => n1339);
   U1383 : AOI221_X1 port map( B1 => n1179, B2 => n3661, C1 => n1180, C2 => 
                           n3693, A => n1344, ZN => n1343);
   U1384 : OAI22_X1 port map( A1 => n1000, A2 => n1182, B1 => n968, B2 => n1183
                           , ZN => n1344);
   U1385 : AOI221_X1 port map( B1 => n1184, B2 => n3725, C1 => n1185, C2 => 
                           n3757, A => n1345, ZN => n1342);
   U1386 : OAI22_X1 port map( A1 => n872, A2 => n1187, B1 => n840, B2 => n1188,
                           ZN => n1345);
   U1387 : AOI221_X1 port map( B1 => n1189, B2 => n3789, C1 => n1190, C2 => 
                           n3821, A => n1346, ZN => n1341);
   U1388 : OAI22_X1 port map( A1 => n680, A2 => n1192, B1 => n648, B2 => n1193,
                           ZN => n1346);
   U1389 : AOI221_X1 port map( B1 => n1194, B2 => n3853, C1 => n1195, C2 => 
                           n3885, A => n1347, ZN => n1340);
   U1390 : OAI22_X1 port map( A1 => n552, A2 => n1197, B1 => n520, B2 => n1198,
                           ZN => n1347);
   U1391 : NAND4_X1 port map( A1 => n1348, A2 => n1349, A3 => n1350, A4 => 
                           n1351, ZN => n1338);
   U1392 : AOI221_X1 port map( B1 => n1203, B2 => n3917, C1 => n1204, C2 => 
                           n3949, A => n1352, ZN => n1351);
   U1393 : OAI22_X1 port map( A1 => n424, A2 => n1206, B1 => n392, B2 => n1207,
                           ZN => n1352);
   U1394 : AOI221_X1 port map( B1 => n1208, B2 => n3981, C1 => n1209, C2 => 
                           n4013, A => n1353, ZN => n1350);
   U1395 : OAI22_X1 port map( A1 => n296, A2 => n1211, B1 => n264, B2 => n1212,
                           ZN => n1353);
   U1396 : AOI221_X1 port map( B1 => n1213, B2 => n143, C1 => n1214, C2 => n15,
                           A => n1354, ZN => n1349);
   U1397 : OAI22_X1 port map( A1 => n79, A2 => n1216, B1 => n207, B2 => n1217, 
                           ZN => n1354);
   U1398 : AOI221_X1 port map( B1 => n1218, B2 => n144, C1 => n1219, C2 => n16,
                           A => n1355, ZN => n1348);
   U1399 : OAI22_X1 port map( A1 => n80, A2 => n1221, B1 => n208, B2 => n1222, 
                           ZN => n1355);
   U1400 : OAI22_X1 port map( A1 => n3628, A2 => n1170, B1 => n1356, B2 => 
                           n1172, ZN => n2582);
   U1401 : NOR2_X1 port map( A1 => n1357, A2 => n1358, ZN => n1356);
   U1402 : NAND4_X1 port map( A1 => n1359, A2 => n1360, A3 => n1361, A4 => 
                           n1362, ZN => n1358);
   U1403 : AOI221_X1 port map( B1 => n1179, B2 => n3660, C1 => n1180, C2 => 
                           n3692, A => n1363, ZN => n1362);
   U1404 : OAI22_X1 port map( A1 => n1001, A2 => n1182, B1 => n969, B2 => n1183
                           , ZN => n1363);
   U1405 : AOI221_X1 port map( B1 => n1184, B2 => n3724, C1 => n1185, C2 => 
                           n3756, A => n1364, ZN => n1361);
   U1406 : OAI22_X1 port map( A1 => n873, A2 => n1187, B1 => n841, B2 => n1188,
                           ZN => n1364);
   U1407 : AOI221_X1 port map( B1 => n1189, B2 => n3788, C1 => n1190, C2 => 
                           n3820, A => n1365, ZN => n1360);
   U1408 : OAI22_X1 port map( A1 => n681, A2 => n1192, B1 => n649, B2 => n1193,
                           ZN => n1365);
   U1409 : AOI221_X1 port map( B1 => n1194, B2 => n3852, C1 => n1195, C2 => 
                           n3884, A => n1366, ZN => n1359);
   U1410 : OAI22_X1 port map( A1 => n553, A2 => n1197, B1 => n521, B2 => n1198,
                           ZN => n1366);
   U1411 : NAND4_X1 port map( A1 => n1367, A2 => n1368, A3 => n1369, A4 => 
                           n1370, ZN => n1357);
   U1412 : AOI221_X1 port map( B1 => n1203, B2 => n3916, C1 => n1204, C2 => 
                           n3948, A => n1371, ZN => n1370);
   U1413 : OAI22_X1 port map( A1 => n425, A2 => n1206, B1 => n393, B2 => n1207,
                           ZN => n1371);
   U1414 : AOI221_X1 port map( B1 => n1208, B2 => n3980, C1 => n1209, C2 => 
                           n4012, A => n1372, ZN => n1369);
   U1415 : OAI22_X1 port map( A1 => n297, A2 => n1211, B1 => n265, B2 => n1212,
                           ZN => n1372);
   U1416 : AOI221_X1 port map( B1 => n1213, B2 => n145, C1 => n1214, C2 => n17,
                           A => n1373, ZN => n1368);
   U1417 : OAI22_X1 port map( A1 => n81, A2 => n1216, B1 => n209, B2 => n1217, 
                           ZN => n1373);
   U1418 : AOI221_X1 port map( B1 => n1218, B2 => n146, C1 => n1219, C2 => n18,
                           A => n1374, ZN => n1367);
   U1419 : OAI22_X1 port map( A1 => n82, A2 => n1221, B1 => n210, B2 => n1222, 
                           ZN => n1374);
   U1420 : OAI22_X1 port map( A1 => n3627, A2 => n1170, B1 => n1375, B2 => 
                           n1172, ZN => n2581);
   U1421 : NOR2_X1 port map( A1 => n1376, A2 => n1377, ZN => n1375);
   U1422 : NAND4_X1 port map( A1 => n1378, A2 => n1379, A3 => n1380, A4 => 
                           n1381, ZN => n1377);
   U1423 : AOI221_X1 port map( B1 => n1179, B2 => n3659, C1 => n1180, C2 => 
                           n3691, A => n1382, ZN => n1381);
   U1424 : OAI22_X1 port map( A1 => n1002, A2 => n1182, B1 => n970, B2 => n1183
                           , ZN => n1382);
   U1425 : AOI221_X1 port map( B1 => n1184, B2 => n3723, C1 => n1185, C2 => 
                           n3755, A => n1383, ZN => n1380);
   U1426 : OAI22_X1 port map( A1 => n874, A2 => n1187, B1 => n842, B2 => n1188,
                           ZN => n1383);
   U1427 : AOI221_X1 port map( B1 => n1189, B2 => n3787, C1 => n1190, C2 => 
                           n3819, A => n1384, ZN => n1379);
   U1428 : OAI22_X1 port map( A1 => n682, A2 => n1192, B1 => n650, B2 => n1193,
                           ZN => n1384);
   U1429 : AOI221_X1 port map( B1 => n1194, B2 => n3851, C1 => n1195, C2 => 
                           n3883, A => n1385, ZN => n1378);
   U1430 : OAI22_X1 port map( A1 => n554, A2 => n1197, B1 => n522, B2 => n1198,
                           ZN => n1385);
   U1431 : NAND4_X1 port map( A1 => n1386, A2 => n1387, A3 => n1388, A4 => 
                           n1389, ZN => n1376);
   U1432 : AOI221_X1 port map( B1 => n1203, B2 => n3915, C1 => n1204, C2 => 
                           n3947, A => n1390, ZN => n1389);
   U1433 : OAI22_X1 port map( A1 => n426, A2 => n1206, B1 => n394, B2 => n1207,
                           ZN => n1390);
   U1434 : AOI221_X1 port map( B1 => n1208, B2 => n3979, C1 => n1209, C2 => 
                           n4011, A => n1391, ZN => n1388);
   U1435 : OAI22_X1 port map( A1 => n298, A2 => n1211, B1 => n266, B2 => n1212,
                           ZN => n1391);
   U1436 : AOI221_X1 port map( B1 => n1213, B2 => n147, C1 => n1214, C2 => n19,
                           A => n1392, ZN => n1387);
   U1437 : OAI22_X1 port map( A1 => n83, A2 => n1216, B1 => n211, B2 => n1217, 
                           ZN => n1392);
   U1438 : AOI221_X1 port map( B1 => n1218, B2 => n148, C1 => n1219, C2 => n20,
                           A => n1393, ZN => n1386);
   U1439 : OAI22_X1 port map( A1 => n84, A2 => n1221, B1 => n212, B2 => n1222, 
                           ZN => n1393);
   U1440 : OAI22_X1 port map( A1 => n3626, A2 => n1170, B1 => n1394, B2 => 
                           n1172, ZN => n2580);
   U1441 : NOR2_X1 port map( A1 => n1395, A2 => n1396, ZN => n1394);
   U1442 : NAND4_X1 port map( A1 => n1397, A2 => n1398, A3 => n1399, A4 => 
                           n1400, ZN => n1396);
   U1443 : AOI221_X1 port map( B1 => n1179, B2 => n3658, C1 => n1180, C2 => 
                           n3690, A => n1401, ZN => n1400);
   U1444 : OAI22_X1 port map( A1 => n1003, A2 => n1182, B1 => n971, B2 => n1183
                           , ZN => n1401);
   U1445 : AOI221_X1 port map( B1 => n1184, B2 => n3722, C1 => n1185, C2 => 
                           n3754, A => n1402, ZN => n1399);
   U1446 : OAI22_X1 port map( A1 => n875, A2 => n1187, B1 => n843, B2 => n1188,
                           ZN => n1402);
   U1447 : AOI221_X1 port map( B1 => n1189, B2 => n3786, C1 => n1190, C2 => 
                           n3818, A => n1403, ZN => n1398);
   U1448 : OAI22_X1 port map( A1 => n683, A2 => n1192, B1 => n651, B2 => n1193,
                           ZN => n1403);
   U1449 : AOI221_X1 port map( B1 => n1194, B2 => n3850, C1 => n1195, C2 => 
                           n3882, A => n1404, ZN => n1397);
   U1450 : OAI22_X1 port map( A1 => n555, A2 => n1197, B1 => n523, B2 => n1198,
                           ZN => n1404);
   U1451 : NAND4_X1 port map( A1 => n1405, A2 => n1406, A3 => n1407, A4 => 
                           n1408, ZN => n1395);
   U1452 : AOI221_X1 port map( B1 => n1203, B2 => n3914, C1 => n1204, C2 => 
                           n3946, A => n1409, ZN => n1408);
   U1453 : OAI22_X1 port map( A1 => n427, A2 => n1206, B1 => n395, B2 => n1207,
                           ZN => n1409);
   U1454 : AOI221_X1 port map( B1 => n1208, B2 => n3978, C1 => n1209, C2 => 
                           n4010, A => n1410, ZN => n1407);
   U1455 : OAI22_X1 port map( A1 => n299, A2 => n1211, B1 => n267, B2 => n1212,
                           ZN => n1410);
   U1456 : AOI221_X1 port map( B1 => n1213, B2 => n149, C1 => n1214, C2 => n21,
                           A => n1411, ZN => n1406);
   U1457 : OAI22_X1 port map( A1 => n85, A2 => n1216, B1 => n213, B2 => n1217, 
                           ZN => n1411);
   U1458 : AOI221_X1 port map( B1 => n1218, B2 => n150, C1 => n1219, C2 => n22,
                           A => n1412, ZN => n1405);
   U1459 : OAI22_X1 port map( A1 => n86, A2 => n1221, B1 => n214, B2 => n1222, 
                           ZN => n1412);
   U1460 : OAI22_X1 port map( A1 => n3625, A2 => n1170, B1 => n1413, B2 => 
                           n1172, ZN => n2579);
   U1461 : NOR2_X1 port map( A1 => n1414, A2 => n1415, ZN => n1413);
   U1462 : NAND4_X1 port map( A1 => n1416, A2 => n1417, A3 => n1418, A4 => 
                           n1419, ZN => n1415);
   U1463 : AOI221_X1 port map( B1 => n1179, B2 => n3657, C1 => n1180, C2 => 
                           n3689, A => n1420, ZN => n1419);
   U1464 : OAI22_X1 port map( A1 => n1004, A2 => n1182, B1 => n972, B2 => n1183
                           , ZN => n1420);
   U1465 : AOI221_X1 port map( B1 => n1184, B2 => n3721, C1 => n1185, C2 => 
                           n3753, A => n1421, ZN => n1418);
   U1466 : OAI22_X1 port map( A1 => n876, A2 => n1187, B1 => n844, B2 => n1188,
                           ZN => n1421);
   U1467 : AOI221_X1 port map( B1 => n1189, B2 => n3785, C1 => n1190, C2 => 
                           n3817, A => n1422, ZN => n1417);
   U1468 : OAI22_X1 port map( A1 => n684, A2 => n1192, B1 => n652, B2 => n1193,
                           ZN => n1422);
   U1469 : AOI221_X1 port map( B1 => n1194, B2 => n3849, C1 => n1195, C2 => 
                           n3881, A => n1423, ZN => n1416);
   U1470 : OAI22_X1 port map( A1 => n556, A2 => n1197, B1 => n524, B2 => n1198,
                           ZN => n1423);
   U1471 : NAND4_X1 port map( A1 => n1424, A2 => n1425, A3 => n1426, A4 => 
                           n1427, ZN => n1414);
   U1472 : AOI221_X1 port map( B1 => n1203, B2 => n3913, C1 => n1204, C2 => 
                           n3945, A => n1428, ZN => n1427);
   U1473 : OAI22_X1 port map( A1 => n428, A2 => n1206, B1 => n396, B2 => n1207,
                           ZN => n1428);
   U1474 : AOI221_X1 port map( B1 => n1208, B2 => n3977, C1 => n1209, C2 => 
                           n4009, A => n1429, ZN => n1426);
   U1475 : OAI22_X1 port map( A1 => n300, A2 => n1211, B1 => n268, B2 => n1212,
                           ZN => n1429);
   U1476 : AOI221_X1 port map( B1 => n1213, B2 => n151, C1 => n1214, C2 => n23,
                           A => n1430, ZN => n1425);
   U1477 : OAI22_X1 port map( A1 => n87, A2 => n1216, B1 => n215, B2 => n1217, 
                           ZN => n1430);
   U1478 : AOI221_X1 port map( B1 => n1218, B2 => n152, C1 => n1219, C2 => n24,
                           A => n1431, ZN => n1424);
   U1479 : OAI22_X1 port map( A1 => n88, A2 => n1221, B1 => n216, B2 => n1222, 
                           ZN => n1431);
   U1480 : OAI22_X1 port map( A1 => n3624, A2 => n1170, B1 => n1432, B2 => 
                           n1172, ZN => n2578);
   U1481 : NOR2_X1 port map( A1 => n1433, A2 => n1434, ZN => n1432);
   U1482 : NAND4_X1 port map( A1 => n1435, A2 => n1436, A3 => n1437, A4 => 
                           n1438, ZN => n1434);
   U1483 : AOI221_X1 port map( B1 => n1179, B2 => n3656, C1 => n1180, C2 => 
                           n3688, A => n1439, ZN => n1438);
   U1484 : OAI22_X1 port map( A1 => n1005, A2 => n1182, B1 => n973, B2 => n1183
                           , ZN => n1439);
   U1485 : AOI221_X1 port map( B1 => n1184, B2 => n3720, C1 => n1185, C2 => 
                           n3752, A => n1440, ZN => n1437);
   U1486 : OAI22_X1 port map( A1 => n877, A2 => n1187, B1 => n845, B2 => n1188,
                           ZN => n1440);
   U1487 : AOI221_X1 port map( B1 => n1189, B2 => n3784, C1 => n1190, C2 => 
                           n3816, A => n1441, ZN => n1436);
   U1488 : OAI22_X1 port map( A1 => n685, A2 => n1192, B1 => n653, B2 => n1193,
                           ZN => n1441);
   U1489 : AOI221_X1 port map( B1 => n1194, B2 => n3848, C1 => n1195, C2 => 
                           n3880, A => n1442, ZN => n1435);
   U1490 : OAI22_X1 port map( A1 => n557, A2 => n1197, B1 => n525, B2 => n1198,
                           ZN => n1442);
   U1491 : NAND4_X1 port map( A1 => n1443, A2 => n1444, A3 => n1445, A4 => 
                           n1446, ZN => n1433);
   U1492 : AOI221_X1 port map( B1 => n1203, B2 => n3912, C1 => n1204, C2 => 
                           n3944, A => n1447, ZN => n1446);
   U1493 : OAI22_X1 port map( A1 => n429, A2 => n1206, B1 => n397, B2 => n1207,
                           ZN => n1447);
   U1494 : AOI221_X1 port map( B1 => n1208, B2 => n3976, C1 => n1209, C2 => 
                           n4008, A => n1448, ZN => n1445);
   U1495 : OAI22_X1 port map( A1 => n301, A2 => n1211, B1 => n269, B2 => n1212,
                           ZN => n1448);
   U1496 : AOI221_X1 port map( B1 => n1213, B2 => n153, C1 => n1214, C2 => n25,
                           A => n1449, ZN => n1444);
   U1497 : OAI22_X1 port map( A1 => n89, A2 => n1216, B1 => n217, B2 => n1217, 
                           ZN => n1449);
   U1498 : AOI221_X1 port map( B1 => n1218, B2 => n154, C1 => n1219, C2 => n26,
                           A => n1450, ZN => n1443);
   U1499 : OAI22_X1 port map( A1 => n90, A2 => n1221, B1 => n218, B2 => n1222, 
                           ZN => n1450);
   U1500 : OAI22_X1 port map( A1 => n3623, A2 => n1170, B1 => n1451, B2 => 
                           n1172, ZN => n2577);
   U1501 : NOR2_X1 port map( A1 => n1452, A2 => n1453, ZN => n1451);
   U1502 : NAND4_X1 port map( A1 => n1454, A2 => n1455, A3 => n1456, A4 => 
                           n1457, ZN => n1453);
   U1503 : AOI221_X1 port map( B1 => n1179, B2 => n3655, C1 => n1180, C2 => 
                           n3687, A => n1458, ZN => n1457);
   U1504 : OAI22_X1 port map( A1 => n1006, A2 => n1182, B1 => n974, B2 => n1183
                           , ZN => n1458);
   U1505 : AOI221_X1 port map( B1 => n1184, B2 => n3719, C1 => n1185, C2 => 
                           n3751, A => n1459, ZN => n1456);
   U1506 : OAI22_X1 port map( A1 => n878, A2 => n1187, B1 => n846, B2 => n1188,
                           ZN => n1459);
   U1507 : AOI221_X1 port map( B1 => n1189, B2 => n3783, C1 => n1190, C2 => 
                           n3815, A => n1460, ZN => n1455);
   U1508 : OAI22_X1 port map( A1 => n686, A2 => n1192, B1 => n654, B2 => n1193,
                           ZN => n1460);
   U1509 : AOI221_X1 port map( B1 => n1194, B2 => n3847, C1 => n1195, C2 => 
                           n3879, A => n1461, ZN => n1454);
   U1510 : OAI22_X1 port map( A1 => n558, A2 => n1197, B1 => n526, B2 => n1198,
                           ZN => n1461);
   U1511 : NAND4_X1 port map( A1 => n1462, A2 => n1463, A3 => n1464, A4 => 
                           n1465, ZN => n1452);
   U1512 : AOI221_X1 port map( B1 => n1203, B2 => n3911, C1 => n1204, C2 => 
                           n3943, A => n1466, ZN => n1465);
   U1513 : OAI22_X1 port map( A1 => n430, A2 => n1206, B1 => n398, B2 => n1207,
                           ZN => n1466);
   U1514 : AOI221_X1 port map( B1 => n1208, B2 => n3975, C1 => n1209, C2 => 
                           n4007, A => n1467, ZN => n1464);
   U1515 : OAI22_X1 port map( A1 => n302, A2 => n1211, B1 => n270, B2 => n1212,
                           ZN => n1467);
   U1516 : AOI221_X1 port map( B1 => n1213, B2 => n155, C1 => n1214, C2 => n27,
                           A => n1468, ZN => n1463);
   U1517 : OAI22_X1 port map( A1 => n91, A2 => n1216, B1 => n219, B2 => n1217, 
                           ZN => n1468);
   U1518 : AOI221_X1 port map( B1 => n1218, B2 => n156, C1 => n1219, C2 => n28,
                           A => n1469, ZN => n1462);
   U1519 : OAI22_X1 port map( A1 => n92, A2 => n1221, B1 => n220, B2 => n1222, 
                           ZN => n1469);
   U1520 : OAI22_X1 port map( A1 => n3622, A2 => n1170, B1 => n1470, B2 => 
                           n1172, ZN => n2576);
   U1521 : NOR2_X1 port map( A1 => n1471, A2 => n1472, ZN => n1470);
   U1522 : NAND4_X1 port map( A1 => n1473, A2 => n1474, A3 => n1475, A4 => 
                           n1476, ZN => n1472);
   U1523 : AOI221_X1 port map( B1 => n1179, B2 => n3654, C1 => n1180, C2 => 
                           n3686, A => n1477, ZN => n1476);
   U1524 : OAI22_X1 port map( A1 => n1007, A2 => n1182, B1 => n975, B2 => n1183
                           , ZN => n1477);
   U1525 : AOI221_X1 port map( B1 => n1184, B2 => n3718, C1 => n1185, C2 => 
                           n3750, A => n1478, ZN => n1475);
   U1526 : OAI22_X1 port map( A1 => n879, A2 => n1187, B1 => n847, B2 => n1188,
                           ZN => n1478);
   U1527 : AOI221_X1 port map( B1 => n1189, B2 => n3782, C1 => n1190, C2 => 
                           n3814, A => n1479, ZN => n1474);
   U1528 : OAI22_X1 port map( A1 => n687, A2 => n1192, B1 => n655, B2 => n1193,
                           ZN => n1479);
   U1529 : AOI221_X1 port map( B1 => n1194, B2 => n3846, C1 => n1195, C2 => 
                           n3878, A => n1480, ZN => n1473);
   U1530 : OAI22_X1 port map( A1 => n559, A2 => n1197, B1 => n527, B2 => n1198,
                           ZN => n1480);
   U1531 : NAND4_X1 port map( A1 => n1481, A2 => n1482, A3 => n1483, A4 => 
                           n1484, ZN => n1471);
   U1532 : AOI221_X1 port map( B1 => n1203, B2 => n3910, C1 => n1204, C2 => 
                           n3942, A => n1485, ZN => n1484);
   U1533 : OAI22_X1 port map( A1 => n431, A2 => n1206, B1 => n399, B2 => n1207,
                           ZN => n1485);
   U1534 : AOI221_X1 port map( B1 => n1208, B2 => n3974, C1 => n1209, C2 => 
                           n4006, A => n1486, ZN => n1483);
   U1535 : OAI22_X1 port map( A1 => n303, A2 => n1211, B1 => n271, B2 => n1212,
                           ZN => n1486);
   U1536 : AOI221_X1 port map( B1 => n1213, B2 => n157, C1 => n1214, C2 => n29,
                           A => n1487, ZN => n1482);
   U1537 : OAI22_X1 port map( A1 => n93, A2 => n1216, B1 => n221, B2 => n1217, 
                           ZN => n1487);
   U1538 : AOI221_X1 port map( B1 => n1218, B2 => n158, C1 => n1219, C2 => n30,
                           A => n1488, ZN => n1481);
   U1539 : OAI22_X1 port map( A1 => n94, A2 => n1221, B1 => n222, B2 => n1222, 
                           ZN => n1488);
   U1540 : OAI22_X1 port map( A1 => n3621, A2 => n1170, B1 => n1489, B2 => 
                           n1172, ZN => n2575);
   U1541 : NOR2_X1 port map( A1 => n1490, A2 => n1491, ZN => n1489);
   U1542 : NAND4_X1 port map( A1 => n1492, A2 => n1493, A3 => n1494, A4 => 
                           n1495, ZN => n1491);
   U1543 : AOI221_X1 port map( B1 => n1179, B2 => n3653, C1 => n1180, C2 => 
                           n3685, A => n1496, ZN => n1495);
   U1544 : OAI22_X1 port map( A1 => n1008, A2 => n1182, B1 => n976, B2 => n1183
                           , ZN => n1496);
   U1545 : AOI221_X1 port map( B1 => n1184, B2 => n3717, C1 => n1185, C2 => 
                           n3749, A => n1497, ZN => n1494);
   U1546 : OAI22_X1 port map( A1 => n880, A2 => n1187, B1 => n848, B2 => n1188,
                           ZN => n1497);
   U1547 : AOI221_X1 port map( B1 => n1189, B2 => n3781, C1 => n1190, C2 => 
                           n3813, A => n1498, ZN => n1493);
   U1548 : OAI22_X1 port map( A1 => n688, A2 => n1192, B1 => n656, B2 => n1193,
                           ZN => n1498);
   U1549 : AOI221_X1 port map( B1 => n1194, B2 => n3845, C1 => n1195, C2 => 
                           n3877, A => n1499, ZN => n1492);
   U1550 : OAI22_X1 port map( A1 => n560, A2 => n1197, B1 => n528, B2 => n1198,
                           ZN => n1499);
   U1551 : NAND4_X1 port map( A1 => n1500, A2 => n1501, A3 => n1502, A4 => 
                           n1503, ZN => n1490);
   U1552 : AOI221_X1 port map( B1 => n1203, B2 => n3909, C1 => n1204, C2 => 
                           n3941, A => n1504, ZN => n1503);
   U1553 : OAI22_X1 port map( A1 => n432, A2 => n1206, B1 => n400, B2 => n1207,
                           ZN => n1504);
   U1554 : AOI221_X1 port map( B1 => n1208, B2 => n3973, C1 => n1209, C2 => 
                           n4005, A => n1505, ZN => n1502);
   U1555 : OAI22_X1 port map( A1 => n304, A2 => n1211, B1 => n272, B2 => n1212,
                           ZN => n1505);
   U1556 : AOI221_X1 port map( B1 => n1213, B2 => n159, C1 => n1214, C2 => n31,
                           A => n1506, ZN => n1501);
   U1557 : OAI22_X1 port map( A1 => n95, A2 => n1216, B1 => n223, B2 => n1217, 
                           ZN => n1506);
   U1558 : AOI221_X1 port map( B1 => n1218, B2 => n160, C1 => n1219, C2 => n32,
                           A => n1507, ZN => n1500);
   U1559 : OAI22_X1 port map( A1 => n96, A2 => n1221, B1 => n224, B2 => n1222, 
                           ZN => n1507);
   U1560 : OAI22_X1 port map( A1 => n3620, A2 => n1170, B1 => n1508, B2 => 
                           n1172, ZN => n2574);
   U1561 : NOR2_X1 port map( A1 => n1509, A2 => n1510, ZN => n1508);
   U1562 : NAND4_X1 port map( A1 => n1511, A2 => n1512, A3 => n1513, A4 => 
                           n1514, ZN => n1510);
   U1563 : AOI221_X1 port map( B1 => n1179, B2 => n3652, C1 => n1180, C2 => 
                           n3684, A => n1515, ZN => n1514);
   U1564 : OAI22_X1 port map( A1 => n1009, A2 => n1182, B1 => n977, B2 => n1183
                           , ZN => n1515);
   U1565 : AOI221_X1 port map( B1 => n1184, B2 => n3716, C1 => n1185, C2 => 
                           n3748, A => n1516, ZN => n1513);
   U1566 : OAI22_X1 port map( A1 => n881, A2 => n1187, B1 => n849, B2 => n1188,
                           ZN => n1516);
   U1567 : AOI221_X1 port map( B1 => n1189, B2 => n3780, C1 => n1190, C2 => 
                           n3812, A => n1517, ZN => n1512);
   U1568 : OAI22_X1 port map( A1 => n689, A2 => n1192, B1 => n657, B2 => n1193,
                           ZN => n1517);
   U1569 : AOI221_X1 port map( B1 => n1194, B2 => n3844, C1 => n1195, C2 => 
                           n3876, A => n1518, ZN => n1511);
   U1570 : OAI22_X1 port map( A1 => n561, A2 => n1197, B1 => n529, B2 => n1198,
                           ZN => n1518);
   U1571 : NAND4_X1 port map( A1 => n1519, A2 => n1520, A3 => n1521, A4 => 
                           n1522, ZN => n1509);
   U1572 : AOI221_X1 port map( B1 => n1203, B2 => n3908, C1 => n1204, C2 => 
                           n3940, A => n1523, ZN => n1522);
   U1573 : OAI22_X1 port map( A1 => n433, A2 => n1206, B1 => n401, B2 => n1207,
                           ZN => n1523);
   U1574 : AOI221_X1 port map( B1 => n1208, B2 => n3972, C1 => n1209, C2 => 
                           n4004, A => n1524, ZN => n1521);
   U1575 : OAI22_X1 port map( A1 => n305, A2 => n1211, B1 => n273, B2 => n1212,
                           ZN => n1524);
   U1576 : AOI221_X1 port map( B1 => n1213, B2 => n161, C1 => n1214, C2 => n33,
                           A => n1525, ZN => n1520);
   U1577 : OAI22_X1 port map( A1 => n97, A2 => n1216, B1 => n225, B2 => n1217, 
                           ZN => n1525);
   U1578 : AOI221_X1 port map( B1 => n1218, B2 => n162, C1 => n1219, C2 => n34,
                           A => n1526, ZN => n1519);
   U1579 : OAI22_X1 port map( A1 => n98, A2 => n1221, B1 => n226, B2 => n1222, 
                           ZN => n1526);
   U1580 : OAI22_X1 port map( A1 => n3619, A2 => n1170, B1 => n1527, B2 => 
                           n1172, ZN => n2573);
   U1581 : NOR2_X1 port map( A1 => n1528, A2 => n1529, ZN => n1527);
   U1582 : NAND4_X1 port map( A1 => n1530, A2 => n1531, A3 => n1532, A4 => 
                           n1533, ZN => n1529);
   U1583 : AOI221_X1 port map( B1 => n1179, B2 => n3651, C1 => n1180, C2 => 
                           n3683, A => n1534, ZN => n1533);
   U1584 : OAI22_X1 port map( A1 => n1010, A2 => n1182, B1 => n978, B2 => n1183
                           , ZN => n1534);
   U1585 : AOI221_X1 port map( B1 => n1184, B2 => n3715, C1 => n1185, C2 => 
                           n3747, A => n1535, ZN => n1532);
   U1586 : OAI22_X1 port map( A1 => n882, A2 => n1187, B1 => n850, B2 => n1188,
                           ZN => n1535);
   U1587 : AOI221_X1 port map( B1 => n1189, B2 => n3779, C1 => n1190, C2 => 
                           n3811, A => n1536, ZN => n1531);
   U1588 : OAI22_X1 port map( A1 => n690, A2 => n1192, B1 => n658, B2 => n1193,
                           ZN => n1536);
   U1589 : AOI221_X1 port map( B1 => n1194, B2 => n3843, C1 => n1195, C2 => 
                           n3875, A => n1537, ZN => n1530);
   U1590 : OAI22_X1 port map( A1 => n562, A2 => n1197, B1 => n530, B2 => n1198,
                           ZN => n1537);
   U1591 : NAND4_X1 port map( A1 => n1538, A2 => n1539, A3 => n1540, A4 => 
                           n1541, ZN => n1528);
   U1592 : AOI221_X1 port map( B1 => n1203, B2 => n3907, C1 => n1204, C2 => 
                           n3939, A => n1542, ZN => n1541);
   U1593 : OAI22_X1 port map( A1 => n434, A2 => n1206, B1 => n402, B2 => n1207,
                           ZN => n1542);
   U1594 : AOI221_X1 port map( B1 => n1208, B2 => n3971, C1 => n1209, C2 => 
                           n4003, A => n1543, ZN => n1540);
   U1595 : OAI22_X1 port map( A1 => n306, A2 => n1211, B1 => n274, B2 => n1212,
                           ZN => n1543);
   U1596 : AOI221_X1 port map( B1 => n1213, B2 => n163, C1 => n1214, C2 => n35,
                           A => n1544, ZN => n1539);
   U1597 : OAI22_X1 port map( A1 => n99, A2 => n1216, B1 => n227, B2 => n1217, 
                           ZN => n1544);
   U1598 : AOI221_X1 port map( B1 => n1218, B2 => n164, C1 => n1219, C2 => n36,
                           A => n1545, ZN => n1538);
   U1599 : OAI22_X1 port map( A1 => n100, A2 => n1221, B1 => n228, B2 => n1222,
                           ZN => n1545);
   U1600 : OAI22_X1 port map( A1 => n3618, A2 => n1170, B1 => n1546, B2 => 
                           n1172, ZN => n2572);
   U1601 : NOR2_X1 port map( A1 => n1547, A2 => n1548, ZN => n1546);
   U1602 : NAND4_X1 port map( A1 => n1549, A2 => n1550, A3 => n1551, A4 => 
                           n1552, ZN => n1548);
   U1603 : AOI221_X1 port map( B1 => n1179, B2 => n3650, C1 => n1180, C2 => 
                           n3682, A => n1553, ZN => n1552);
   U1604 : OAI22_X1 port map( A1 => n1011, A2 => n1182, B1 => n979, B2 => n1183
                           , ZN => n1553);
   U1605 : AOI221_X1 port map( B1 => n1184, B2 => n3714, C1 => n1185, C2 => 
                           n3746, A => n1554, ZN => n1551);
   U1606 : OAI22_X1 port map( A1 => n883, A2 => n1187, B1 => n851, B2 => n1188,
                           ZN => n1554);
   U1607 : AOI221_X1 port map( B1 => n1189, B2 => n3778, C1 => n1190, C2 => 
                           n3810, A => n1555, ZN => n1550);
   U1608 : OAI22_X1 port map( A1 => n691, A2 => n1192, B1 => n659, B2 => n1193,
                           ZN => n1555);
   U1609 : AOI221_X1 port map( B1 => n1194, B2 => n3842, C1 => n1195, C2 => 
                           n3874, A => n1556, ZN => n1549);
   U1610 : OAI22_X1 port map( A1 => n563, A2 => n1197, B1 => n531, B2 => n1198,
                           ZN => n1556);
   U1611 : NAND4_X1 port map( A1 => n1557, A2 => n1558, A3 => n1559, A4 => 
                           n1560, ZN => n1547);
   U1612 : AOI221_X1 port map( B1 => n1203, B2 => n3906, C1 => n1204, C2 => 
                           n3938, A => n1561, ZN => n1560);
   U1613 : OAI22_X1 port map( A1 => n435, A2 => n1206, B1 => n403, B2 => n1207,
                           ZN => n1561);
   U1614 : AOI221_X1 port map( B1 => n1208, B2 => n3970, C1 => n1209, C2 => 
                           n4002, A => n1562, ZN => n1559);
   U1615 : OAI22_X1 port map( A1 => n307, A2 => n1211, B1 => n275, B2 => n1212,
                           ZN => n1562);
   U1616 : AOI221_X1 port map( B1 => n1213, B2 => n165, C1 => n1214, C2 => n37,
                           A => n1563, ZN => n1558);
   U1617 : OAI22_X1 port map( A1 => n101, A2 => n1216, B1 => n229, B2 => n1217,
                           ZN => n1563);
   U1618 : AOI221_X1 port map( B1 => n1218, B2 => n166, C1 => n1219, C2 => n38,
                           A => n1564, ZN => n1557);
   U1619 : OAI22_X1 port map( A1 => n102, A2 => n1221, B1 => n230, B2 => n1222,
                           ZN => n1564);
   U1620 : OAI22_X1 port map( A1 => n3617, A2 => n1170, B1 => n1565, B2 => 
                           n1172, ZN => n2571);
   U1621 : NOR2_X1 port map( A1 => n1566, A2 => n1567, ZN => n1565);
   U1622 : NAND4_X1 port map( A1 => n1568, A2 => n1569, A3 => n1570, A4 => 
                           n1571, ZN => n1567);
   U1623 : AOI221_X1 port map( B1 => n1179, B2 => n3649, C1 => n1180, C2 => 
                           n3681, A => n1572, ZN => n1571);
   U1624 : OAI22_X1 port map( A1 => n1012, A2 => n1182, B1 => n980, B2 => n1183
                           , ZN => n1572);
   U1625 : AOI221_X1 port map( B1 => n1184, B2 => n3713, C1 => n1185, C2 => 
                           n3745, A => n1573, ZN => n1570);
   U1626 : OAI22_X1 port map( A1 => n884, A2 => n1187, B1 => n852, B2 => n1188,
                           ZN => n1573);
   U1627 : AOI221_X1 port map( B1 => n1189, B2 => n3777, C1 => n1190, C2 => 
                           n3809, A => n1574, ZN => n1569);
   U1628 : OAI22_X1 port map( A1 => n692, A2 => n1192, B1 => n660, B2 => n1193,
                           ZN => n1574);
   U1629 : AOI221_X1 port map( B1 => n1194, B2 => n3841, C1 => n1195, C2 => 
                           n3873, A => n1575, ZN => n1568);
   U1630 : OAI22_X1 port map( A1 => n564, A2 => n1197, B1 => n532, B2 => n1198,
                           ZN => n1575);
   U1631 : NAND4_X1 port map( A1 => n1576, A2 => n1577, A3 => n1578, A4 => 
                           n1579, ZN => n1566);
   U1632 : AOI221_X1 port map( B1 => n1203, B2 => n3905, C1 => n1204, C2 => 
                           n3937, A => n1580, ZN => n1579);
   U1633 : OAI22_X1 port map( A1 => n436, A2 => n1206, B1 => n404, B2 => n1207,
                           ZN => n1580);
   U1634 : AOI221_X1 port map( B1 => n1208, B2 => n3969, C1 => n1209, C2 => 
                           n4001, A => n1581, ZN => n1578);
   U1635 : OAI22_X1 port map( A1 => n308, A2 => n1211, B1 => n276, B2 => n1212,
                           ZN => n1581);
   U1636 : AOI221_X1 port map( B1 => n1213, B2 => n167, C1 => n1214, C2 => n39,
                           A => n1582, ZN => n1577);
   U1637 : OAI22_X1 port map( A1 => n103, A2 => n1216, B1 => n231, B2 => n1217,
                           ZN => n1582);
   U1638 : AOI221_X1 port map( B1 => n1218, B2 => n168, C1 => n1219, C2 => n40,
                           A => n1583, ZN => n1576);
   U1639 : OAI22_X1 port map( A1 => n104, A2 => n1221, B1 => n232, B2 => n1222,
                           ZN => n1583);
   U1640 : OAI22_X1 port map( A1 => n3616, A2 => n1170, B1 => n1584, B2 => 
                           n1172, ZN => n2570);
   U1641 : NOR2_X1 port map( A1 => n1585, A2 => n1586, ZN => n1584);
   U1642 : NAND4_X1 port map( A1 => n1587, A2 => n1588, A3 => n1589, A4 => 
                           n1590, ZN => n1586);
   U1643 : AOI221_X1 port map( B1 => n1179, B2 => n3648, C1 => n1180, C2 => 
                           n3680, A => n1591, ZN => n1590);
   U1644 : OAI22_X1 port map( A1 => n1013, A2 => n1182, B1 => n981, B2 => n1183
                           , ZN => n1591);
   U1645 : AOI221_X1 port map( B1 => n1184, B2 => n3712, C1 => n1185, C2 => 
                           n3744, A => n1592, ZN => n1589);
   U1646 : OAI22_X1 port map( A1 => n885, A2 => n1187, B1 => n853, B2 => n1188,
                           ZN => n1592);
   U1647 : AOI221_X1 port map( B1 => n1189, B2 => n3776, C1 => n1190, C2 => 
                           n3808, A => n1593, ZN => n1588);
   U1648 : OAI22_X1 port map( A1 => n693, A2 => n1192, B1 => n661, B2 => n1193,
                           ZN => n1593);
   U1649 : AOI221_X1 port map( B1 => n1194, B2 => n3840, C1 => n1195, C2 => 
                           n3872, A => n1594, ZN => n1587);
   U1650 : OAI22_X1 port map( A1 => n565, A2 => n1197, B1 => n533, B2 => n1198,
                           ZN => n1594);
   U1651 : NAND4_X1 port map( A1 => n1595, A2 => n1596, A3 => n1597, A4 => 
                           n1598, ZN => n1585);
   U1652 : AOI221_X1 port map( B1 => n1203, B2 => n3904, C1 => n1204, C2 => 
                           n3936, A => n1599, ZN => n1598);
   U1653 : OAI22_X1 port map( A1 => n437, A2 => n1206, B1 => n405, B2 => n1207,
                           ZN => n1599);
   U1654 : AOI221_X1 port map( B1 => n1208, B2 => n3968, C1 => n1209, C2 => 
                           n4000, A => n1600, ZN => n1597);
   U1655 : OAI22_X1 port map( A1 => n309, A2 => n1211, B1 => n277, B2 => n1212,
                           ZN => n1600);
   U1656 : AOI221_X1 port map( B1 => n1213, B2 => n169, C1 => n1214, C2 => n41,
                           A => n1601, ZN => n1596);
   U1657 : OAI22_X1 port map( A1 => n105, A2 => n1216, B1 => n233, B2 => n1217,
                           ZN => n1601);
   U1658 : AOI221_X1 port map( B1 => n1218, B2 => n170, C1 => n1219, C2 => n42,
                           A => n1602, ZN => n1595);
   U1659 : OAI22_X1 port map( A1 => n106, A2 => n1221, B1 => n234, B2 => n1222,
                           ZN => n1602);
   U1660 : OAI22_X1 port map( A1 => n3615, A2 => n1170, B1 => n1603, B2 => 
                           n1172, ZN => n2569);
   U1661 : NOR2_X1 port map( A1 => n1604, A2 => n1605, ZN => n1603);
   U1662 : NAND4_X1 port map( A1 => n1606, A2 => n1607, A3 => n1608, A4 => 
                           n1609, ZN => n1605);
   U1663 : AOI221_X1 port map( B1 => n1179, B2 => n3647, C1 => n1180, C2 => 
                           n3679, A => n1610, ZN => n1609);
   U1664 : OAI22_X1 port map( A1 => n1014, A2 => n1182, B1 => n982, B2 => n1183
                           , ZN => n1610);
   U1665 : AOI221_X1 port map( B1 => n1184, B2 => n3711, C1 => n1185, C2 => 
                           n3743, A => n1611, ZN => n1608);
   U1666 : OAI22_X1 port map( A1 => n886, A2 => n1187, B1 => n854, B2 => n1188,
                           ZN => n1611);
   U1667 : AOI221_X1 port map( B1 => n1189, B2 => n3775, C1 => n1190, C2 => 
                           n3807, A => n1612, ZN => n1607);
   U1668 : OAI22_X1 port map( A1 => n694, A2 => n1192, B1 => n662, B2 => n1193,
                           ZN => n1612);
   U1669 : AOI221_X1 port map( B1 => n1194, B2 => n3839, C1 => n1195, C2 => 
                           n3871, A => n1613, ZN => n1606);
   U1670 : OAI22_X1 port map( A1 => n566, A2 => n1197, B1 => n534, B2 => n1198,
                           ZN => n1613);
   U1671 : NAND4_X1 port map( A1 => n1614, A2 => n1615, A3 => n1616, A4 => 
                           n1617, ZN => n1604);
   U1672 : AOI221_X1 port map( B1 => n1203, B2 => n3903, C1 => n1204, C2 => 
                           n3935, A => n1618, ZN => n1617);
   U1673 : OAI22_X1 port map( A1 => n438, A2 => n1206, B1 => n406, B2 => n1207,
                           ZN => n1618);
   U1674 : AOI221_X1 port map( B1 => n1208, B2 => n3967, C1 => n1209, C2 => 
                           n3999, A => n1619, ZN => n1616);
   U1675 : OAI22_X1 port map( A1 => n310, A2 => n1211, B1 => n278, B2 => n1212,
                           ZN => n1619);
   U1676 : AOI221_X1 port map( B1 => n1213, B2 => n171, C1 => n1214, C2 => n43,
                           A => n1620, ZN => n1615);
   U1677 : OAI22_X1 port map( A1 => n107, A2 => n1216, B1 => n235, B2 => n1217,
                           ZN => n1620);
   U1678 : AOI221_X1 port map( B1 => n1218, B2 => n172, C1 => n1219, C2 => n44,
                           A => n1621, ZN => n1614);
   U1679 : OAI22_X1 port map( A1 => n108, A2 => n1221, B1 => n236, B2 => n1222,
                           ZN => n1621);
   U1680 : OAI22_X1 port map( A1 => n2526, A2 => n1170, B1 => n1622, B2 => 
                           n1172, ZN => n2568);
   U1681 : NOR2_X1 port map( A1 => n1623, A2 => n1624, ZN => n1622);
   U1682 : NAND4_X1 port map( A1 => n1625, A2 => n1626, A3 => n1627, A4 => 
                           n1628, ZN => n1624);
   U1683 : AOI221_X1 port map( B1 => n1179, B2 => n3646, C1 => n1180, C2 => 
                           n3678, A => n1629, ZN => n1628);
   U1684 : OAI22_X1 port map( A1 => n1015, A2 => n1182, B1 => n983, B2 => n1183
                           , ZN => n1629);
   U1685 : AOI221_X1 port map( B1 => n1184, B2 => n3710, C1 => n1185, C2 => 
                           n3742, A => n1630, ZN => n1627);
   U1686 : OAI22_X1 port map( A1 => n887, A2 => n1187, B1 => n855, B2 => n1188,
                           ZN => n1630);
   U1687 : AOI221_X1 port map( B1 => n1189, B2 => n3774, C1 => n1190, C2 => 
                           n3806, A => n1631, ZN => n1626);
   U1688 : OAI22_X1 port map( A1 => n695, A2 => n1192, B1 => n663, B2 => n1193,
                           ZN => n1631);
   U1689 : AOI221_X1 port map( B1 => n1194, B2 => n3838, C1 => n1195, C2 => 
                           n3870, A => n1632, ZN => n1625);
   U1690 : OAI22_X1 port map( A1 => n567, A2 => n1197, B1 => n535, B2 => n1198,
                           ZN => n1632);
   U1691 : NAND4_X1 port map( A1 => n1633, A2 => n1634, A3 => n1635, A4 => 
                           n1636, ZN => n1623);
   U1692 : AOI221_X1 port map( B1 => n1203, B2 => n3902, C1 => n1204, C2 => 
                           n3934, A => n1637, ZN => n1636);
   U1693 : OAI22_X1 port map( A1 => n439, A2 => n1206, B1 => n407, B2 => n1207,
                           ZN => n1637);
   U1694 : AOI221_X1 port map( B1 => n1208, B2 => n3966, C1 => n1209, C2 => 
                           n3998, A => n1638, ZN => n1635);
   U1695 : OAI22_X1 port map( A1 => n311, A2 => n1211, B1 => n279, B2 => n1212,
                           ZN => n1638);
   U1696 : AOI221_X1 port map( B1 => n1213, B2 => n173, C1 => n1214, C2 => n45,
                           A => n1639, ZN => n1634);
   U1697 : OAI22_X1 port map( A1 => n109, A2 => n1216, B1 => n237, B2 => n1217,
                           ZN => n1639);
   U1698 : AOI221_X1 port map( B1 => n1218, B2 => n174, C1 => n1219, C2 => n46,
                           A => n1640, ZN => n1633);
   U1699 : OAI22_X1 port map( A1 => n110, A2 => n1221, B1 => n238, B2 => n1222,
                           ZN => n1640);
   U1700 : OAI22_X1 port map( A1 => n2525, A2 => n1170, B1 => n1641, B2 => 
                           n1172, ZN => n2567);
   U1701 : NOR2_X1 port map( A1 => n1642, A2 => n1643, ZN => n1641);
   U1702 : NAND4_X1 port map( A1 => n1644, A2 => n1645, A3 => n1646, A4 => 
                           n1647, ZN => n1643);
   U1703 : AOI221_X1 port map( B1 => n1179, B2 => n3645, C1 => n1180, C2 => 
                           n3677, A => n1648, ZN => n1647);
   U1704 : OAI22_X1 port map( A1 => n1016, A2 => n1182, B1 => n984, B2 => n1183
                           , ZN => n1648);
   U1705 : AOI221_X1 port map( B1 => n1184, B2 => n3709, C1 => n1185, C2 => 
                           n3741, A => n1649, ZN => n1646);
   U1706 : OAI22_X1 port map( A1 => n888, A2 => n1187, B1 => n856, B2 => n1188,
                           ZN => n1649);
   U1707 : AOI221_X1 port map( B1 => n1189, B2 => n3773, C1 => n1190, C2 => 
                           n3805, A => n1650, ZN => n1645);
   U1708 : OAI22_X1 port map( A1 => n696, A2 => n1192, B1 => n664, B2 => n1193,
                           ZN => n1650);
   U1709 : AOI221_X1 port map( B1 => n1194, B2 => n3837, C1 => n1195, C2 => 
                           n3869, A => n1651, ZN => n1644);
   U1710 : OAI22_X1 port map( A1 => n568, A2 => n1197, B1 => n536, B2 => n1198,
                           ZN => n1651);
   U1711 : NAND4_X1 port map( A1 => n1652, A2 => n1653, A3 => n1654, A4 => 
                           n1655, ZN => n1642);
   U1712 : AOI221_X1 port map( B1 => n1203, B2 => n3901, C1 => n1204, C2 => 
                           n3933, A => n1656, ZN => n1655);
   U1713 : OAI22_X1 port map( A1 => n440, A2 => n1206, B1 => n408, B2 => n1207,
                           ZN => n1656);
   U1714 : AOI221_X1 port map( B1 => n1208, B2 => n3965, C1 => n1209, C2 => 
                           n3997, A => n1657, ZN => n1654);
   U1715 : OAI22_X1 port map( A1 => n312, A2 => n1211, B1 => n280, B2 => n1212,
                           ZN => n1657);
   U1716 : AOI221_X1 port map( B1 => n1213, B2 => n175, C1 => n1214, C2 => n47,
                           A => n1658, ZN => n1653);
   U1717 : OAI22_X1 port map( A1 => n111, A2 => n1216, B1 => n239, B2 => n1217,
                           ZN => n1658);
   U1718 : AOI221_X1 port map( B1 => n1218, B2 => n176, C1 => n1219, C2 => n48,
                           A => n1659, ZN => n1652);
   U1719 : OAI22_X1 port map( A1 => n112, A2 => n1221, B1 => n240, B2 => n1222,
                           ZN => n1659);
   U1720 : OAI22_X1 port map( A1 => n2524, A2 => n1170, B1 => n1660, B2 => 
                           n1172, ZN => n2566);
   U1721 : NOR2_X1 port map( A1 => n1661, A2 => n1662, ZN => n1660);
   U1722 : NAND4_X1 port map( A1 => n1663, A2 => n1664, A3 => n1665, A4 => 
                           n1666, ZN => n1662);
   U1723 : AOI221_X1 port map( B1 => n1179, B2 => n3644, C1 => n1180, C2 => 
                           n3676, A => n1667, ZN => n1666);
   U1724 : OAI22_X1 port map( A1 => n1017, A2 => n1182, B1 => n985, B2 => n1183
                           , ZN => n1667);
   U1725 : AOI221_X1 port map( B1 => n1184, B2 => n3708, C1 => n1185, C2 => 
                           n3740, A => n1668, ZN => n1665);
   U1726 : OAI22_X1 port map( A1 => n889, A2 => n1187, B1 => n857, B2 => n1188,
                           ZN => n1668);
   U1727 : AOI221_X1 port map( B1 => n1189, B2 => n3772, C1 => n1190, C2 => 
                           n3804, A => n1669, ZN => n1664);
   U1728 : OAI22_X1 port map( A1 => n697, A2 => n1192, B1 => n665, B2 => n1193,
                           ZN => n1669);
   U1729 : AOI221_X1 port map( B1 => n1194, B2 => n3836, C1 => n1195, C2 => 
                           n3868, A => n1670, ZN => n1663);
   U1730 : OAI22_X1 port map( A1 => n569, A2 => n1197, B1 => n537, B2 => n1198,
                           ZN => n1670);
   U1731 : NAND4_X1 port map( A1 => n1671, A2 => n1672, A3 => n1673, A4 => 
                           n1674, ZN => n1661);
   U1732 : AOI221_X1 port map( B1 => n1203, B2 => n3900, C1 => n1204, C2 => 
                           n3932, A => n1675, ZN => n1674);
   U1733 : OAI22_X1 port map( A1 => n441, A2 => n1206, B1 => n409, B2 => n1207,
                           ZN => n1675);
   U1734 : AOI221_X1 port map( B1 => n1208, B2 => n3964, C1 => n1209, C2 => 
                           n3996, A => n1676, ZN => n1673);
   U1735 : OAI22_X1 port map( A1 => n313, A2 => n1211, B1 => n281, B2 => n1212,
                           ZN => n1676);
   U1736 : AOI221_X1 port map( B1 => n1213, B2 => n177, C1 => n1214, C2 => n49,
                           A => n1677, ZN => n1672);
   U1737 : OAI22_X1 port map( A1 => n113, A2 => n1216, B1 => n241, B2 => n1217,
                           ZN => n1677);
   U1738 : AOI221_X1 port map( B1 => n1218, B2 => n178, C1 => n1219, C2 => n50,
                           A => n1678, ZN => n1671);
   U1739 : OAI22_X1 port map( A1 => n114, A2 => n1221, B1 => n242, B2 => n1222,
                           ZN => n1678);
   U1740 : OAI22_X1 port map( A1 => n2523, A2 => n1170, B1 => n1679, B2 => 
                           n1172, ZN => n2565);
   U1741 : NOR2_X1 port map( A1 => n1680, A2 => n1681, ZN => n1679);
   U1742 : NAND4_X1 port map( A1 => n1682, A2 => n1683, A3 => n1684, A4 => 
                           n1685, ZN => n1681);
   U1743 : AOI221_X1 port map( B1 => n1179, B2 => n3643, C1 => n1180, C2 => 
                           n3675, A => n1686, ZN => n1685);
   U1744 : OAI22_X1 port map( A1 => n1018, A2 => n1182, B1 => n986, B2 => n1183
                           , ZN => n1686);
   U1745 : AOI221_X1 port map( B1 => n1184, B2 => n3707, C1 => n1185, C2 => 
                           n3739, A => n1687, ZN => n1684);
   U1746 : OAI22_X1 port map( A1 => n890, A2 => n1187, B1 => n858, B2 => n1188,
                           ZN => n1687);
   U1747 : AOI221_X1 port map( B1 => n1189, B2 => n3771, C1 => n1190, C2 => 
                           n3803, A => n1688, ZN => n1683);
   U1748 : OAI22_X1 port map( A1 => n698, A2 => n1192, B1 => n666, B2 => n1193,
                           ZN => n1688);
   U1749 : AOI221_X1 port map( B1 => n1194, B2 => n3835, C1 => n1195, C2 => 
                           n3867, A => n1689, ZN => n1682);
   U1750 : OAI22_X1 port map( A1 => n570, A2 => n1197, B1 => n538, B2 => n1198,
                           ZN => n1689);
   U1751 : NAND4_X1 port map( A1 => n1690, A2 => n1691, A3 => n1692, A4 => 
                           n1693, ZN => n1680);
   U1752 : AOI221_X1 port map( B1 => n1203, B2 => n3899, C1 => n1204, C2 => 
                           n3931, A => n1694, ZN => n1693);
   U1753 : OAI22_X1 port map( A1 => n442, A2 => n1206, B1 => n410, B2 => n1207,
                           ZN => n1694);
   U1754 : AOI221_X1 port map( B1 => n1208, B2 => n3963, C1 => n1209, C2 => 
                           n3995, A => n1695, ZN => n1692);
   U1755 : OAI22_X1 port map( A1 => n314, A2 => n1211, B1 => n282, B2 => n1212,
                           ZN => n1695);
   U1756 : AOI221_X1 port map( B1 => n1213, B2 => n179, C1 => n1214, C2 => n51,
                           A => n1696, ZN => n1691);
   U1757 : OAI22_X1 port map( A1 => n115, A2 => n1216, B1 => n243, B2 => n1217,
                           ZN => n1696);
   U1758 : AOI221_X1 port map( B1 => n1218, B2 => n180, C1 => n1219, C2 => n52,
                           A => n1697, ZN => n1690);
   U1759 : OAI22_X1 port map( A1 => n116, A2 => n1221, B1 => n244, B2 => n1222,
                           ZN => n1697);
   U1760 : OAI22_X1 port map( A1 => n2522, A2 => n1170, B1 => n1698, B2 => 
                           n1172, ZN => n2564);
   U1761 : NOR2_X1 port map( A1 => n1699, A2 => n1700, ZN => n1698);
   U1762 : NAND4_X1 port map( A1 => n1701, A2 => n1702, A3 => n1703, A4 => 
                           n1704, ZN => n1700);
   U1763 : AOI221_X1 port map( B1 => n1179, B2 => n3642, C1 => n1180, C2 => 
                           n3674, A => n1705, ZN => n1704);
   U1764 : OAI22_X1 port map( A1 => n1019, A2 => n1182, B1 => n987, B2 => n1183
                           , ZN => n1705);
   U1765 : AOI221_X1 port map( B1 => n1184, B2 => n3706, C1 => n1185, C2 => 
                           n3738, A => n1706, ZN => n1703);
   U1766 : OAI22_X1 port map( A1 => n891, A2 => n1187, B1 => n859, B2 => n1188,
                           ZN => n1706);
   U1767 : AOI221_X1 port map( B1 => n1189, B2 => n3770, C1 => n1190, C2 => 
                           n3802, A => n1707, ZN => n1702);
   U1768 : OAI22_X1 port map( A1 => n699, A2 => n1192, B1 => n667, B2 => n1193,
                           ZN => n1707);
   U1769 : AOI221_X1 port map( B1 => n1194, B2 => n3834, C1 => n1195, C2 => 
                           n3866, A => n1708, ZN => n1701);
   U1770 : OAI22_X1 port map( A1 => n571, A2 => n1197, B1 => n539, B2 => n1198,
                           ZN => n1708);
   U1771 : NAND4_X1 port map( A1 => n1709, A2 => n1710, A3 => n1711, A4 => 
                           n1712, ZN => n1699);
   U1772 : AOI221_X1 port map( B1 => n1203, B2 => n3898, C1 => n1204, C2 => 
                           n3930, A => n1713, ZN => n1712);
   U1773 : OAI22_X1 port map( A1 => n443, A2 => n1206, B1 => n411, B2 => n1207,
                           ZN => n1713);
   U1774 : AOI221_X1 port map( B1 => n1208, B2 => n3962, C1 => n1209, C2 => 
                           n3994, A => n1714, ZN => n1711);
   U1775 : OAI22_X1 port map( A1 => n315, A2 => n1211, B1 => n283, B2 => n1212,
                           ZN => n1714);
   U1776 : AOI221_X1 port map( B1 => n1213, B2 => n181, C1 => n1214, C2 => n53,
                           A => n1715, ZN => n1710);
   U1777 : OAI22_X1 port map( A1 => n117, A2 => n1216, B1 => n245, B2 => n1217,
                           ZN => n1715);
   U1778 : AOI221_X1 port map( B1 => n1218, B2 => n182, C1 => n1219, C2 => n54,
                           A => n1716, ZN => n1709);
   U1779 : OAI22_X1 port map( A1 => n118, A2 => n1221, B1 => n246, B2 => n1222,
                           ZN => n1716);
   U1780 : OAI22_X1 port map( A1 => n2521, A2 => n1170, B1 => n1717, B2 => 
                           n1172, ZN => n2563);
   U1781 : NOR2_X1 port map( A1 => n1718, A2 => n1719, ZN => n1717);
   U1782 : NAND4_X1 port map( A1 => n1720, A2 => n1721, A3 => n1722, A4 => 
                           n1723, ZN => n1719);
   U1783 : AOI221_X1 port map( B1 => n1179, B2 => n3641, C1 => n1180, C2 => 
                           n3673, A => n1724, ZN => n1723);
   U1784 : OAI22_X1 port map( A1 => n1020, A2 => n1182, B1 => n988, B2 => n1183
                           , ZN => n1724);
   U1785 : AOI221_X1 port map( B1 => n1184, B2 => n3705, C1 => n1185, C2 => 
                           n3737, A => n1725, ZN => n1722);
   U1786 : OAI22_X1 port map( A1 => n892, A2 => n1187, B1 => n860, B2 => n1188,
                           ZN => n1725);
   U1787 : AOI221_X1 port map( B1 => n1189, B2 => n3769, C1 => n1190, C2 => 
                           n3801, A => n1726, ZN => n1721);
   U1788 : OAI22_X1 port map( A1 => n700, A2 => n1192, B1 => n668, B2 => n1193,
                           ZN => n1726);
   U1789 : AOI221_X1 port map( B1 => n1194, B2 => n3833, C1 => n1195, C2 => 
                           n3865, A => n1727, ZN => n1720);
   U1790 : OAI22_X1 port map( A1 => n572, A2 => n1197, B1 => n540, B2 => n1198,
                           ZN => n1727);
   U1791 : NAND4_X1 port map( A1 => n1728, A2 => n1729, A3 => n1730, A4 => 
                           n1731, ZN => n1718);
   U1792 : AOI221_X1 port map( B1 => n1203, B2 => n3897, C1 => n1204, C2 => 
                           n3929, A => n1732, ZN => n1731);
   U1793 : OAI22_X1 port map( A1 => n444, A2 => n1206, B1 => n412, B2 => n1207,
                           ZN => n1732);
   U1794 : AOI221_X1 port map( B1 => n1208, B2 => n3961, C1 => n1209, C2 => 
                           n3993, A => n1733, ZN => n1730);
   U1795 : OAI22_X1 port map( A1 => n316, A2 => n1211, B1 => n284, B2 => n1212,
                           ZN => n1733);
   U1796 : AOI221_X1 port map( B1 => n1213, B2 => n183, C1 => n1214, C2 => n55,
                           A => n1734, ZN => n1729);
   U1797 : OAI22_X1 port map( A1 => n119, A2 => n1216, B1 => n247, B2 => n1217,
                           ZN => n1734);
   U1798 : AOI221_X1 port map( B1 => n1218, B2 => n184, C1 => n1219, C2 => n56,
                           A => n1735, ZN => n1728);
   U1799 : OAI22_X1 port map( A1 => n120, A2 => n1221, B1 => n248, B2 => n1222,
                           ZN => n1735);
   U1800 : OAI22_X1 port map( A1 => n2520, A2 => n1170, B1 => n1736, B2 => 
                           n1172, ZN => n2562);
   U1801 : NOR2_X1 port map( A1 => n1737, A2 => n1738, ZN => n1736);
   U1802 : NAND4_X1 port map( A1 => n1739, A2 => n1740, A3 => n1741, A4 => 
                           n1742, ZN => n1738);
   U1803 : AOI221_X1 port map( B1 => n1179, B2 => n3640, C1 => n1180, C2 => 
                           n3672, A => n1743, ZN => n1742);
   U1804 : OAI22_X1 port map( A1 => n1021, A2 => n1182, B1 => n989, B2 => n1183
                           , ZN => n1743);
   U1805 : AOI221_X1 port map( B1 => n1184, B2 => n3704, C1 => n1185, C2 => 
                           n3736, A => n1744, ZN => n1741);
   U1806 : OAI22_X1 port map( A1 => n893, A2 => n1187, B1 => n861, B2 => n1188,
                           ZN => n1744);
   U1807 : AOI221_X1 port map( B1 => n1189, B2 => n3768, C1 => n1190, C2 => 
                           n3800, A => n1745, ZN => n1740);
   U1808 : OAI22_X1 port map( A1 => n701, A2 => n1192, B1 => n669, B2 => n1193,
                           ZN => n1745);
   U1809 : AOI221_X1 port map( B1 => n1194, B2 => n3832, C1 => n1195, C2 => 
                           n3864, A => n1746, ZN => n1739);
   U1810 : OAI22_X1 port map( A1 => n573, A2 => n1197, B1 => n541, B2 => n1198,
                           ZN => n1746);
   U1811 : NAND4_X1 port map( A1 => n1747, A2 => n1748, A3 => n1749, A4 => 
                           n1750, ZN => n1737);
   U1812 : AOI221_X1 port map( B1 => n1203, B2 => n3896, C1 => n1204, C2 => 
                           n3928, A => n1751, ZN => n1750);
   U1813 : OAI22_X1 port map( A1 => n445, A2 => n1206, B1 => n413, B2 => n1207,
                           ZN => n1751);
   U1814 : AOI221_X1 port map( B1 => n1208, B2 => n3960, C1 => n1209, C2 => 
                           n3992, A => n1752, ZN => n1749);
   U1815 : OAI22_X1 port map( A1 => n317, A2 => n1211, B1 => n285, B2 => n1212,
                           ZN => n1752);
   U1816 : AOI221_X1 port map( B1 => n1213, B2 => n185, C1 => n1214, C2 => n57,
                           A => n1753, ZN => n1748);
   U1817 : OAI22_X1 port map( A1 => n121, A2 => n1216, B1 => n249, B2 => n1217,
                           ZN => n1753);
   U1818 : AOI221_X1 port map( B1 => n1218, B2 => n186, C1 => n1219, C2 => n58,
                           A => n1754, ZN => n1747);
   U1819 : OAI22_X1 port map( A1 => n122, A2 => n1221, B1 => n250, B2 => n1222,
                           ZN => n1754);
   U1820 : OAI22_X1 port map( A1 => n2519, A2 => n1170, B1 => n1755, B2 => 
                           n1172, ZN => n2561);
   U1821 : NOR2_X1 port map( A1 => n1756, A2 => n1757, ZN => n1755);
   U1822 : NAND4_X1 port map( A1 => n1758, A2 => n1759, A3 => n1760, A4 => 
                           n1761, ZN => n1757);
   U1823 : AOI221_X1 port map( B1 => n1179, B2 => n3639, C1 => n1180, C2 => 
                           n3671, A => n1762, ZN => n1761);
   U1824 : OAI22_X1 port map( A1 => n1022, A2 => n1182, B1 => n990, B2 => n1183
                           , ZN => n1762);
   U1825 : AOI221_X1 port map( B1 => n1184, B2 => n3703, C1 => n1185, C2 => 
                           n3735, A => n1763, ZN => n1760);
   U1826 : OAI22_X1 port map( A1 => n894, A2 => n1187, B1 => n862, B2 => n1188,
                           ZN => n1763);
   U1827 : AOI221_X1 port map( B1 => n1189, B2 => n3767, C1 => n1190, C2 => 
                           n3799, A => n1764, ZN => n1759);
   U1828 : OAI22_X1 port map( A1 => n702, A2 => n1192, B1 => n670, B2 => n1193,
                           ZN => n1764);
   U1829 : AOI221_X1 port map( B1 => n1194, B2 => n3831, C1 => n1195, C2 => 
                           n3863, A => n1765, ZN => n1758);
   U1830 : OAI22_X1 port map( A1 => n574, A2 => n1197, B1 => n542, B2 => n1198,
                           ZN => n1765);
   U1831 : NAND4_X1 port map( A1 => n1766, A2 => n1767, A3 => n1768, A4 => 
                           n1769, ZN => n1756);
   U1832 : AOI221_X1 port map( B1 => n1203, B2 => n3895, C1 => n1204, C2 => 
                           n3927, A => n1770, ZN => n1769);
   U1833 : OAI22_X1 port map( A1 => n446, A2 => n1206, B1 => n414, B2 => n1207,
                           ZN => n1770);
   U1834 : AOI221_X1 port map( B1 => n1208, B2 => n3959, C1 => n1209, C2 => 
                           n3991, A => n1771, ZN => n1768);
   U1835 : OAI22_X1 port map( A1 => n318, A2 => n1211, B1 => n286, B2 => n1212,
                           ZN => n1771);
   U1836 : AOI221_X1 port map( B1 => n1213, B2 => n187, C1 => n1214, C2 => n59,
                           A => n1772, ZN => n1767);
   U1837 : OAI22_X1 port map( A1 => n123, A2 => n1216, B1 => n251, B2 => n1217,
                           ZN => n1772);
   U1838 : AOI221_X1 port map( B1 => n1218, B2 => n188, C1 => n1219, C2 => n60,
                           A => n1773, ZN => n1766);
   U1839 : OAI22_X1 port map( A1 => n124, A2 => n1221, B1 => n252, B2 => n1222,
                           ZN => n1773);
   U1840 : OAI22_X1 port map( A1 => n2518, A2 => n1170, B1 => n1774, B2 => 
                           n1172, ZN => n2560);
   U1841 : NOR2_X1 port map( A1 => n1775, A2 => n1776, ZN => n1774);
   U1842 : NAND4_X1 port map( A1 => n1777, A2 => n1778, A3 => n1779, A4 => 
                           n1780, ZN => n1776);
   U1843 : AOI221_X1 port map( B1 => n1179, B2 => n3638, C1 => n1180, C2 => 
                           n3670, A => n1781, ZN => n1780);
   U1844 : OAI22_X1 port map( A1 => n1023, A2 => n1182, B1 => n991, B2 => n1183
                           , ZN => n1781);
   U1845 : AOI221_X1 port map( B1 => n1184, B2 => n3702, C1 => n1185, C2 => 
                           n3734, A => n1782, ZN => n1779);
   U1846 : OAI22_X1 port map( A1 => n895, A2 => n1187, B1 => n863, B2 => n1188,
                           ZN => n1782);
   U1847 : AOI221_X1 port map( B1 => n1189, B2 => n3766, C1 => n1190, C2 => 
                           n3798, A => n1783, ZN => n1778);
   U1848 : OAI22_X1 port map( A1 => n703, A2 => n1192, B1 => n671, B2 => n1193,
                           ZN => n1783);
   U1849 : AOI221_X1 port map( B1 => n1194, B2 => n3830, C1 => n1195, C2 => 
                           n3862, A => n1784, ZN => n1777);
   U1850 : OAI22_X1 port map( A1 => n575, A2 => n1197, B1 => n543, B2 => n1198,
                           ZN => n1784);
   U1851 : NAND4_X1 port map( A1 => n1785, A2 => n1786, A3 => n1787, A4 => 
                           n1788, ZN => n1775);
   U1852 : AOI221_X1 port map( B1 => n1203, B2 => n3894, C1 => n1204, C2 => 
                           n3926, A => n1789, ZN => n1788);
   U1853 : OAI22_X1 port map( A1 => n447, A2 => n1206, B1 => n415, B2 => n1207,
                           ZN => n1789);
   U1854 : AOI221_X1 port map( B1 => n1208, B2 => n3958, C1 => n1209, C2 => 
                           n3990, A => n1790, ZN => n1787);
   U1855 : OAI22_X1 port map( A1 => n319, A2 => n1211, B1 => n287, B2 => n1212,
                           ZN => n1790);
   U1856 : AOI221_X1 port map( B1 => n1213, B2 => n189, C1 => n1214, C2 => n61,
                           A => n1791, ZN => n1786);
   U1857 : OAI22_X1 port map( A1 => n125, A2 => n1216, B1 => n253, B2 => n1217,
                           ZN => n1791);
   U1858 : AOI221_X1 port map( B1 => n1218, B2 => n190, C1 => n1219, C2 => n62,
                           A => n1792, ZN => n1785);
   U1859 : OAI22_X1 port map( A1 => n126, A2 => n1221, B1 => n254, B2 => n1222,
                           ZN => n1792);
   U1860 : OAI22_X1 port map( A1 => n2517, A2 => n1170, B1 => n1793, B2 => 
                           n1172, ZN => n2559);
   U1861 : NOR2_X1 port map( A1 => n1794, A2 => n1795, ZN => n1793);
   U1862 : NAND4_X1 port map( A1 => n1796, A2 => n1797, A3 => n1798, A4 => 
                           n1799, ZN => n1795);
   U1863 : AOI221_X1 port map( B1 => n1179, B2 => n3637, C1 => n1180, C2 => 
                           n3669, A => n1800, ZN => n1799);
   U1864 : OAI22_X1 port map( A1 => n1024, A2 => n1182, B1 => n992, B2 => n1183
                           , ZN => n1800);
   U1865 : AOI221_X1 port map( B1 => n1184, B2 => n3701, C1 => n1185, C2 => 
                           n3733, A => n1805, ZN => n1798);
   U1866 : OAI22_X1 port map( A1 => n896, A2 => n1187, B1 => n864, B2 => n1188,
                           ZN => n1805);
   U1867 : AND3_X1 port map( A1 => ADD_RD1(3), A2 => n1808, A3 => ADD_RD1(4), 
                           ZN => n1801);
   U1868 : AND3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(0), A3 => 
                           ADD_RD1(4), ZN => n1803);
   U1869 : AOI221_X1 port map( B1 => n1189, B2 => n3765, C1 => n1190, C2 => 
                           n3797, A => n1809, ZN => n1797);
   U1870 : OAI22_X1 port map( A1 => n704, A2 => n1192, B1 => n672, B2 => n1193,
                           ZN => n1809);
   U1871 : AOI221_X1 port map( B1 => n1194, B2 => n3829, C1 => n1195, C2 => 
                           n3861, A => n1812, ZN => n1796);
   U1872 : OAI22_X1 port map( A1 => n576, A2 => n1197, B1 => n544, B2 => n1198,
                           ZN => n1812);
   U1873 : AND3_X1 port map( A1 => n1808, A2 => n1813, A3 => ADD_RD1(4), ZN => 
                           n1810);
   U1874 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => n1813, A3 => ADD_RD1(4), 
                           ZN => n1811);
   U1875 : NAND4_X1 port map( A1 => n1814, A2 => n1815, A3 => n1816, A4 => 
                           n1817, ZN => n1794);
   U1876 : AOI221_X1 port map( B1 => n1203, B2 => n3893, C1 => n1204, C2 => 
                           n3925, A => n1818, ZN => n1817);
   U1877 : OAI22_X1 port map( A1 => n448, A2 => n1206, B1 => n416, B2 => n1207,
                           ZN => n1818);
   U1878 : AOI221_X1 port map( B1 => n1208, B2 => n3957, C1 => n1209, C2 => 
                           n3989, A => n1821, ZN => n1816);
   U1879 : OAI22_X1 port map( A1 => n320, A2 => n1211, B1 => n288, B2 => n1212,
                           ZN => n1821);
   U1880 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n1813, 
                           ZN => n1819);
   U1881 : NOR3_X1 port map( A1 => n1808, A2 => ADD_RD1(4), A3 => n1813, ZN => 
                           n1820);
   U1882 : INV_X1 port map( A => ADD_RD1(3), ZN => n1813);
   U1883 : AOI221_X1 port map( B1 => n1213, B2 => n191, C1 => n1214, C2 => n63,
                           A => n1822, ZN => n1815);
   U1884 : OAI22_X1 port map( A1 => n127, A2 => n1216, B1 => n255, B2 => n1217,
                           ZN => n1822);
   U1885 : AND2_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), ZN => n1802);
   U1886 : AND2_X1 port map( A1 => ADD_RD1(2), A2 => n1825, ZN => n1804);
   U1887 : AOI221_X1 port map( B1 => n1218, B2 => n192, C1 => n1219, C2 => n64,
                           A => n1826, ZN => n1814);
   U1888 : OAI22_X1 port map( A1 => n128, A2 => n1221, B1 => n256, B2 => n1222,
                           ZN => n1826);
   U1889 : NOR2_X1 port map( A1 => n1825, A2 => ADD_RD1(2), ZN => n1806);
   U1890 : INV_X1 port map( A => ADD_RD1(1), ZN => n1825);
   U1891 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n1808, 
                           ZN => n1823);
   U1892 : INV_X1 port map( A => ADD_RD1(0), ZN => n1808);
   U1893 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n1807);
   U1894 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n1824);
   U1895 : OAI22_X1 port map( A1 => n2516, A2 => n1828, B1 => n1829, B2 => 
                           n1830, ZN => n2558);
   U1896 : NOR2_X1 port map( A1 => n1831, A2 => n1832, ZN => n1829);
   U1897 : NAND4_X1 port map( A1 => n1833, A2 => n1834, A3 => n1835, A4 => 
                           n1836, ZN => n1832);
   U1898 : AOI221_X1 port map( B1 => n1837, B2 => n3668, C1 => n1838, C2 => 
                           n3700, A => n1839, ZN => n1836);
   U1899 : OAI22_X1 port map( A1 => n993, A2 => n1840, B1 => n961, B2 => n1841,
                           ZN => n1839);
   U1900 : AOI221_X1 port map( B1 => n1842, B2 => n3732, C1 => n1843, C2 => 
                           n3764, A => n1844, ZN => n1835);
   U1901 : OAI22_X1 port map( A1 => n865, A2 => n1845, B1 => n833, B2 => n1846,
                           ZN => n1844);
   U1902 : AOI221_X1 port map( B1 => n1847, B2 => n3796, C1 => n1848, C2 => 
                           n3828, A => n1849, ZN => n1834);
   U1903 : OAI22_X1 port map( A1 => n673, A2 => n1850, B1 => n641, B2 => n1851,
                           ZN => n1849);
   U1904 : AOI221_X1 port map( B1 => n1852, B2 => n3860, C1 => n1853, C2 => 
                           n3892, A => n1854, ZN => n1833);
   U1905 : OAI22_X1 port map( A1 => n545, A2 => n1855, B1 => n513, B2 => n1856,
                           ZN => n1854);
   U1906 : NAND4_X1 port map( A1 => n1857, A2 => n1858, A3 => n1859, A4 => 
                           n1860, ZN => n1831);
   U1907 : AOI221_X1 port map( B1 => n1861, B2 => n3924, C1 => n1862, C2 => 
                           n3956, A => n1863, ZN => n1860);
   U1908 : OAI22_X1 port map( A1 => n417, A2 => n1864, B1 => n385, B2 => n1865,
                           ZN => n1863);
   U1909 : AOI221_X1 port map( B1 => n1866, B2 => n3988, C1 => n1867, C2 => 
                           n4020, A => n1868, ZN => n1859);
   U1910 : OAI22_X1 port map( A1 => n289, A2 => n1869, B1 => n257, B2 => n1870,
                           ZN => n1868);
   U1911 : AOI221_X1 port map( B1 => n1871, B2 => n129, C1 => n1872, C2 => n1, 
                           A => n1873, ZN => n1858);
   U1912 : OAI22_X1 port map( A1 => n65, A2 => n1874, B1 => n193, B2 => n1875, 
                           ZN => n1873);
   U1913 : AOI221_X1 port map( B1 => n1876, B2 => n130, C1 => n1877, C2 => n2, 
                           A => n1878, ZN => n1857);
   U1914 : OAI22_X1 port map( A1 => n66, A2 => n1879, B1 => n194, B2 => n1880, 
                           ZN => n1878);
   U1915 : OAI22_X1 port map( A1 => n2515, A2 => n1828, B1 => n1881, B2 => 
                           n1830, ZN => n2557);
   U1916 : NOR2_X1 port map( A1 => n1882, A2 => n1883, ZN => n1881);
   U1917 : NAND4_X1 port map( A1 => n1884, A2 => n1885, A3 => n1886, A4 => 
                           n1887, ZN => n1883);
   U1918 : AOI221_X1 port map( B1 => n1837, B2 => n3667, C1 => n1838, C2 => 
                           n3699, A => n1888, ZN => n1887);
   U1919 : OAI22_X1 port map( A1 => n994, A2 => n1840, B1 => n962, B2 => n1841,
                           ZN => n1888);
   U1920 : AOI221_X1 port map( B1 => n1842, B2 => n3731, C1 => n1843, C2 => 
                           n3763, A => n1889, ZN => n1886);
   U1921 : OAI22_X1 port map( A1 => n866, A2 => n1845, B1 => n834, B2 => n1846,
                           ZN => n1889);
   U1922 : AOI221_X1 port map( B1 => n1847, B2 => n3795, C1 => n1848, C2 => 
                           n3827, A => n1890, ZN => n1885);
   U1923 : OAI22_X1 port map( A1 => n674, A2 => n1850, B1 => n642, B2 => n1851,
                           ZN => n1890);
   U1924 : AOI221_X1 port map( B1 => n1852, B2 => n3859, C1 => n1853, C2 => 
                           n3891, A => n1891, ZN => n1884);
   U1925 : OAI22_X1 port map( A1 => n546, A2 => n1855, B1 => n514, B2 => n1856,
                           ZN => n1891);
   U1926 : NAND4_X1 port map( A1 => n1892, A2 => n1893, A3 => n1894, A4 => 
                           n1895, ZN => n1882);
   U1927 : AOI221_X1 port map( B1 => n1861, B2 => n3923, C1 => n1862, C2 => 
                           n3955, A => n1896, ZN => n1895);
   U1928 : OAI22_X1 port map( A1 => n418, A2 => n1864, B1 => n386, B2 => n1865,
                           ZN => n1896);
   U1929 : AOI221_X1 port map( B1 => n1866, B2 => n3987, C1 => n1867, C2 => 
                           n4019, A => n1897, ZN => n1894);
   U1930 : OAI22_X1 port map( A1 => n290, A2 => n1869, B1 => n258, B2 => n1870,
                           ZN => n1897);
   U1931 : AOI221_X1 port map( B1 => n1871, B2 => n131, C1 => n1872, C2 => n3, 
                           A => n1898, ZN => n1893);
   U1932 : OAI22_X1 port map( A1 => n67, A2 => n1874, B1 => n195, B2 => n1875, 
                           ZN => n1898);
   U1933 : AOI221_X1 port map( B1 => n1876, B2 => n132, C1 => n1877, C2 => n4, 
                           A => n1899, ZN => n1892);
   U1934 : OAI22_X1 port map( A1 => n68, A2 => n1879, B1 => n196, B2 => n1880, 
                           ZN => n1899);
   U1935 : OAI22_X1 port map( A1 => n2514, A2 => n1828, B1 => n1900, B2 => 
                           n1830, ZN => n2556);
   U1936 : NOR2_X1 port map( A1 => n1901, A2 => n1902, ZN => n1900);
   U1937 : NAND4_X1 port map( A1 => n1903, A2 => n1904, A3 => n1905, A4 => 
                           n1906, ZN => n1902);
   U1938 : AOI221_X1 port map( B1 => n1837, B2 => n3666, C1 => n1838, C2 => 
                           n3698, A => n1907, ZN => n1906);
   U1939 : OAI22_X1 port map( A1 => n995, A2 => n1840, B1 => n963, B2 => n1841,
                           ZN => n1907);
   U1940 : AOI221_X1 port map( B1 => n1842, B2 => n3730, C1 => n1843, C2 => 
                           n3762, A => n1908, ZN => n1905);
   U1941 : OAI22_X1 port map( A1 => n867, A2 => n1845, B1 => n835, B2 => n1846,
                           ZN => n1908);
   U1942 : AOI221_X1 port map( B1 => n1847, B2 => n3794, C1 => n1848, C2 => 
                           n3826, A => n1909, ZN => n1904);
   U1943 : OAI22_X1 port map( A1 => n675, A2 => n1850, B1 => n643, B2 => n1851,
                           ZN => n1909);
   U1944 : AOI221_X1 port map( B1 => n1852, B2 => n3858, C1 => n1853, C2 => 
                           n3890, A => n1910, ZN => n1903);
   U1945 : OAI22_X1 port map( A1 => n547, A2 => n1855, B1 => n515, B2 => n1856,
                           ZN => n1910);
   U1946 : NAND4_X1 port map( A1 => n1911, A2 => n1912, A3 => n1913, A4 => 
                           n1914, ZN => n1901);
   U1947 : AOI221_X1 port map( B1 => n1861, B2 => n3922, C1 => n1862, C2 => 
                           n3954, A => n1915, ZN => n1914);
   U1948 : OAI22_X1 port map( A1 => n419, A2 => n1864, B1 => n387, B2 => n1865,
                           ZN => n1915);
   U1949 : AOI221_X1 port map( B1 => n1866, B2 => n3986, C1 => n1867, C2 => 
                           n4018, A => n1916, ZN => n1913);
   U1950 : OAI22_X1 port map( A1 => n291, A2 => n1869, B1 => n259, B2 => n1870,
                           ZN => n1916);
   U1951 : AOI221_X1 port map( B1 => n1871, B2 => n133, C1 => n1872, C2 => n5, 
                           A => n1917, ZN => n1912);
   U1952 : OAI22_X1 port map( A1 => n69, A2 => n1874, B1 => n197, B2 => n1875, 
                           ZN => n1917);
   U1953 : AOI221_X1 port map( B1 => n1876, B2 => n134, C1 => n1877, C2 => n6, 
                           A => n1918, ZN => n1911);
   U1954 : OAI22_X1 port map( A1 => n70, A2 => n1879, B1 => n198, B2 => n1880, 
                           ZN => n1918);
   U1955 : OAI22_X1 port map( A1 => n2513, A2 => n1828, B1 => n1919, B2 => 
                           n1830, ZN => n2555);
   U1956 : NOR2_X1 port map( A1 => n1920, A2 => n1921, ZN => n1919);
   U1957 : NAND4_X1 port map( A1 => n1922, A2 => n1923, A3 => n1924, A4 => 
                           n1925, ZN => n1921);
   U1958 : AOI221_X1 port map( B1 => n1837, B2 => n3665, C1 => n1838, C2 => 
                           n3697, A => n1926, ZN => n1925);
   U1959 : OAI22_X1 port map( A1 => n996, A2 => n1840, B1 => n964, B2 => n1841,
                           ZN => n1926);
   U1960 : AOI221_X1 port map( B1 => n1842, B2 => n3729, C1 => n1843, C2 => 
                           n3761, A => n1927, ZN => n1924);
   U1961 : OAI22_X1 port map( A1 => n868, A2 => n1845, B1 => n836, B2 => n1846,
                           ZN => n1927);
   U1962 : AOI221_X1 port map( B1 => n1847, B2 => n3793, C1 => n1848, C2 => 
                           n3825, A => n1928, ZN => n1923);
   U1963 : OAI22_X1 port map( A1 => n676, A2 => n1850, B1 => n644, B2 => n1851,
                           ZN => n1928);
   U1964 : AOI221_X1 port map( B1 => n1852, B2 => n3857, C1 => n1853, C2 => 
                           n3889, A => n1929, ZN => n1922);
   U1965 : OAI22_X1 port map( A1 => n548, A2 => n1855, B1 => n516, B2 => n1856,
                           ZN => n1929);
   U1966 : NAND4_X1 port map( A1 => n1930, A2 => n1931, A3 => n1932, A4 => 
                           n1933, ZN => n1920);
   U1967 : AOI221_X1 port map( B1 => n1861, B2 => n3921, C1 => n1862, C2 => 
                           n3953, A => n1934, ZN => n1933);
   U1968 : OAI22_X1 port map( A1 => n420, A2 => n1864, B1 => n388, B2 => n1865,
                           ZN => n1934);
   U1969 : AOI221_X1 port map( B1 => n1866, B2 => n3985, C1 => n1867, C2 => 
                           n4017, A => n1935, ZN => n1932);
   U1970 : OAI22_X1 port map( A1 => n292, A2 => n1869, B1 => n260, B2 => n1870,
                           ZN => n1935);
   U1971 : AOI221_X1 port map( B1 => n1871, B2 => n135, C1 => n1872, C2 => n7, 
                           A => n1936, ZN => n1931);
   U1972 : OAI22_X1 port map( A1 => n71, A2 => n1874, B1 => n199, B2 => n1875, 
                           ZN => n1936);
   U1973 : AOI221_X1 port map( B1 => n1876, B2 => n136, C1 => n1877, C2 => n8, 
                           A => n1937, ZN => n1930);
   U1974 : OAI22_X1 port map( A1 => n72, A2 => n1879, B1 => n200, B2 => n1880, 
                           ZN => n1937);
   U1975 : OAI22_X1 port map( A1 => n2512, A2 => n1828, B1 => n1938, B2 => 
                           n1830, ZN => n2554);
   U1976 : NOR2_X1 port map( A1 => n1939, A2 => n1940, ZN => n1938);
   U1977 : NAND4_X1 port map( A1 => n1941, A2 => n1942, A3 => n1943, A4 => 
                           n1944, ZN => n1940);
   U1978 : AOI221_X1 port map( B1 => n1837, B2 => n3664, C1 => n1838, C2 => 
                           n3696, A => n1945, ZN => n1944);
   U1979 : OAI22_X1 port map( A1 => n997, A2 => n1840, B1 => n965, B2 => n1841,
                           ZN => n1945);
   U1980 : AOI221_X1 port map( B1 => n1842, B2 => n3728, C1 => n1843, C2 => 
                           n3760, A => n1946, ZN => n1943);
   U1981 : OAI22_X1 port map( A1 => n869, A2 => n1845, B1 => n837, B2 => n1846,
                           ZN => n1946);
   U1982 : AOI221_X1 port map( B1 => n1847, B2 => n3792, C1 => n1848, C2 => 
                           n3824, A => n1947, ZN => n1942);
   U1983 : OAI22_X1 port map( A1 => n677, A2 => n1850, B1 => n645, B2 => n1851,
                           ZN => n1947);
   U1984 : AOI221_X1 port map( B1 => n1852, B2 => n3856, C1 => n1853, C2 => 
                           n3888, A => n1948, ZN => n1941);
   U1985 : OAI22_X1 port map( A1 => n549, A2 => n1855, B1 => n517, B2 => n1856,
                           ZN => n1948);
   U1986 : NAND4_X1 port map( A1 => n1949, A2 => n1950, A3 => n1951, A4 => 
                           n1952, ZN => n1939);
   U1987 : AOI221_X1 port map( B1 => n1861, B2 => n3920, C1 => n1862, C2 => 
                           n3952, A => n1953, ZN => n1952);
   U1988 : OAI22_X1 port map( A1 => n421, A2 => n1864, B1 => n389, B2 => n1865,
                           ZN => n1953);
   U1989 : AOI221_X1 port map( B1 => n1866, B2 => n3984, C1 => n1867, C2 => 
                           n4016, A => n1954, ZN => n1951);
   U1990 : OAI22_X1 port map( A1 => n293, A2 => n1869, B1 => n261, B2 => n1870,
                           ZN => n1954);
   U1991 : AOI221_X1 port map( B1 => n1871, B2 => n137, C1 => n1872, C2 => n9, 
                           A => n1955, ZN => n1950);
   U1992 : OAI22_X1 port map( A1 => n73, A2 => n1874, B1 => n201, B2 => n1875, 
                           ZN => n1955);
   U1993 : AOI221_X1 port map( B1 => n1876, B2 => n138, C1 => n1877, C2 => n10,
                           A => n1956, ZN => n1949);
   U1994 : OAI22_X1 port map( A1 => n74, A2 => n1879, B1 => n202, B2 => n1880, 
                           ZN => n1956);
   U1995 : OAI22_X1 port map( A1 => n2511, A2 => n1828, B1 => n1957, B2 => 
                           n1830, ZN => n2553);
   U1996 : NOR2_X1 port map( A1 => n1958, A2 => n1959, ZN => n1957);
   U1997 : NAND4_X1 port map( A1 => n1960, A2 => n1961, A3 => n1962, A4 => 
                           n1963, ZN => n1959);
   U1998 : AOI221_X1 port map( B1 => n1837, B2 => n3663, C1 => n1838, C2 => 
                           n3695, A => n1964, ZN => n1963);
   U1999 : OAI22_X1 port map( A1 => n998, A2 => n1840, B1 => n966, B2 => n1841,
                           ZN => n1964);
   U2000 : AOI221_X1 port map( B1 => n1842, B2 => n3727, C1 => n1843, C2 => 
                           n3759, A => n1965, ZN => n1962);
   U2001 : OAI22_X1 port map( A1 => n870, A2 => n1845, B1 => n838, B2 => n1846,
                           ZN => n1965);
   U2002 : AOI221_X1 port map( B1 => n1847, B2 => n3791, C1 => n1848, C2 => 
                           n3823, A => n1966, ZN => n1961);
   U2003 : OAI22_X1 port map( A1 => n678, A2 => n1850, B1 => n646, B2 => n1851,
                           ZN => n1966);
   U2004 : AOI221_X1 port map( B1 => n1852, B2 => n3855, C1 => n1853, C2 => 
                           n3887, A => n1967, ZN => n1960);
   U2005 : OAI22_X1 port map( A1 => n550, A2 => n1855, B1 => n518, B2 => n1856,
                           ZN => n1967);
   U2006 : NAND4_X1 port map( A1 => n1968, A2 => n1969, A3 => n1970, A4 => 
                           n1971, ZN => n1958);
   U2007 : AOI221_X1 port map( B1 => n1861, B2 => n3919, C1 => n1862, C2 => 
                           n3951, A => n1972, ZN => n1971);
   U2008 : OAI22_X1 port map( A1 => n422, A2 => n1864, B1 => n390, B2 => n1865,
                           ZN => n1972);
   U2009 : AOI221_X1 port map( B1 => n1866, B2 => n3983, C1 => n1867, C2 => 
                           n4015, A => n1973, ZN => n1970);
   U2010 : OAI22_X1 port map( A1 => n294, A2 => n1869, B1 => n262, B2 => n1870,
                           ZN => n1973);
   U2011 : AOI221_X1 port map( B1 => n1871, B2 => n139, C1 => n1872, C2 => n11,
                           A => n1974, ZN => n1969);
   U2012 : OAI22_X1 port map( A1 => n75, A2 => n1874, B1 => n203, B2 => n1875, 
                           ZN => n1974);
   U2013 : AOI221_X1 port map( B1 => n1876, B2 => n140, C1 => n1877, C2 => n12,
                           A => n1975, ZN => n1968);
   U2014 : OAI22_X1 port map( A1 => n76, A2 => n1879, B1 => n204, B2 => n1880, 
                           ZN => n1975);
   U2015 : OAI22_X1 port map( A1 => n2510, A2 => n1828, B1 => n1976, B2 => 
                           n1830, ZN => n2552);
   U2016 : NOR2_X1 port map( A1 => n1977, A2 => n1978, ZN => n1976);
   U2017 : NAND4_X1 port map( A1 => n1979, A2 => n1980, A3 => n1981, A4 => 
                           n1982, ZN => n1978);
   U2018 : AOI221_X1 port map( B1 => n1837, B2 => n3662, C1 => n1838, C2 => 
                           n3694, A => n1983, ZN => n1982);
   U2019 : OAI22_X1 port map( A1 => n999, A2 => n1840, B1 => n967, B2 => n1841,
                           ZN => n1983);
   U2020 : AOI221_X1 port map( B1 => n1842, B2 => n3726, C1 => n1843, C2 => 
                           n3758, A => n1984, ZN => n1981);
   U2021 : OAI22_X1 port map( A1 => n871, A2 => n1845, B1 => n839, B2 => n1846,
                           ZN => n1984);
   U2022 : AOI221_X1 port map( B1 => n1847, B2 => n3790, C1 => n1848, C2 => 
                           n3822, A => n1985, ZN => n1980);
   U2023 : OAI22_X1 port map( A1 => n679, A2 => n1850, B1 => n647, B2 => n1851,
                           ZN => n1985);
   U2024 : AOI221_X1 port map( B1 => n1852, B2 => n3854, C1 => n1853, C2 => 
                           n3886, A => n1986, ZN => n1979);
   U2025 : OAI22_X1 port map( A1 => n551, A2 => n1855, B1 => n519, B2 => n1856,
                           ZN => n1986);
   U2026 : NAND4_X1 port map( A1 => n1987, A2 => n1988, A3 => n1989, A4 => 
                           n1990, ZN => n1977);
   U2027 : AOI221_X1 port map( B1 => n1861, B2 => n3918, C1 => n1862, C2 => 
                           n3950, A => n1991, ZN => n1990);
   U2028 : OAI22_X1 port map( A1 => n423, A2 => n1864, B1 => n391, B2 => n1865,
                           ZN => n1991);
   U2029 : AOI221_X1 port map( B1 => n1866, B2 => n3982, C1 => n1867, C2 => 
                           n4014, A => n1992, ZN => n1989);
   U2030 : OAI22_X1 port map( A1 => n295, A2 => n1869, B1 => n263, B2 => n1870,
                           ZN => n1992);
   U2031 : AOI221_X1 port map( B1 => n1871, B2 => n141, C1 => n1872, C2 => n13,
                           A => n1993, ZN => n1988);
   U2032 : OAI22_X1 port map( A1 => n77, A2 => n1874, B1 => n205, B2 => n1875, 
                           ZN => n1993);
   U2033 : AOI221_X1 port map( B1 => n1876, B2 => n142, C1 => n1877, C2 => n14,
                           A => n1994, ZN => n1987);
   U2034 : OAI22_X1 port map( A1 => n78, A2 => n1879, B1 => n206, B2 => n1880, 
                           ZN => n1994);
   U2035 : OAI22_X1 port map( A1 => n2509, A2 => n1828, B1 => n1995, B2 => 
                           n1830, ZN => n2551);
   U2036 : NOR2_X1 port map( A1 => n1996, A2 => n1997, ZN => n1995);
   U2037 : NAND4_X1 port map( A1 => n1998, A2 => n1999, A3 => n2000, A4 => 
                           n2001, ZN => n1997);
   U2038 : AOI221_X1 port map( B1 => n1837, B2 => n3661, C1 => n1838, C2 => 
                           n3693, A => n2002, ZN => n2001);
   U2039 : OAI22_X1 port map( A1 => n1000, A2 => n1840, B1 => n968, B2 => n1841
                           , ZN => n2002);
   U2040 : AOI221_X1 port map( B1 => n1842, B2 => n3725, C1 => n1843, C2 => 
                           n3757, A => n2003, ZN => n2000);
   U2041 : OAI22_X1 port map( A1 => n872, A2 => n1845, B1 => n840, B2 => n1846,
                           ZN => n2003);
   U2042 : AOI221_X1 port map( B1 => n1847, B2 => n3789, C1 => n1848, C2 => 
                           n3821, A => n2004, ZN => n1999);
   U2043 : OAI22_X1 port map( A1 => n680, A2 => n1850, B1 => n648, B2 => n1851,
                           ZN => n2004);
   U2044 : AOI221_X1 port map( B1 => n1852, B2 => n3853, C1 => n1853, C2 => 
                           n3885, A => n2005, ZN => n1998);
   U2045 : OAI22_X1 port map( A1 => n552, A2 => n1855, B1 => n520, B2 => n1856,
                           ZN => n2005);
   U2046 : NAND4_X1 port map( A1 => n2006, A2 => n2007, A3 => n2008, A4 => 
                           n2009, ZN => n1996);
   U2047 : AOI221_X1 port map( B1 => n1861, B2 => n3917, C1 => n1862, C2 => 
                           n3949, A => n2010, ZN => n2009);
   U2048 : OAI22_X1 port map( A1 => n424, A2 => n1864, B1 => n392, B2 => n1865,
                           ZN => n2010);
   U2049 : AOI221_X1 port map( B1 => n1866, B2 => n3981, C1 => n1867, C2 => 
                           n4013, A => n2011, ZN => n2008);
   U2050 : OAI22_X1 port map( A1 => n296, A2 => n1869, B1 => n264, B2 => n1870,
                           ZN => n2011);
   U2051 : AOI221_X1 port map( B1 => n1871, B2 => n143, C1 => n1872, C2 => n15,
                           A => n2012, ZN => n2007);
   U2052 : OAI22_X1 port map( A1 => n79, A2 => n1874, B1 => n207, B2 => n1875, 
                           ZN => n2012);
   U2053 : AOI221_X1 port map( B1 => n1876, B2 => n144, C1 => n1877, C2 => n16,
                           A => n2013, ZN => n2006);
   U2054 : OAI22_X1 port map( A1 => n80, A2 => n1879, B1 => n208, B2 => n1880, 
                           ZN => n2013);
   U2055 : OAI22_X1 port map( A1 => n2508, A2 => n1828, B1 => n2014, B2 => 
                           n1830, ZN => n2550);
   U2056 : NOR2_X1 port map( A1 => n2015, A2 => n2016, ZN => n2014);
   U2057 : NAND4_X1 port map( A1 => n2017, A2 => n2018, A3 => n2019, A4 => 
                           n2020, ZN => n2016);
   U2058 : AOI221_X1 port map( B1 => n1837, B2 => n3660, C1 => n1838, C2 => 
                           n3692, A => n2021, ZN => n2020);
   U2059 : OAI22_X1 port map( A1 => n1001, A2 => n1840, B1 => n969, B2 => n1841
                           , ZN => n2021);
   U2060 : AOI221_X1 port map( B1 => n1842, B2 => n3724, C1 => n1843, C2 => 
                           n3756, A => n2022, ZN => n2019);
   U2061 : OAI22_X1 port map( A1 => n873, A2 => n1845, B1 => n841, B2 => n1846,
                           ZN => n2022);
   U2062 : AOI221_X1 port map( B1 => n1847, B2 => n3788, C1 => n1848, C2 => 
                           n3820, A => n2023, ZN => n2018);
   U2063 : OAI22_X1 port map( A1 => n681, A2 => n1850, B1 => n649, B2 => n1851,
                           ZN => n2023);
   U2064 : AOI221_X1 port map( B1 => n1852, B2 => n3852, C1 => n1853, C2 => 
                           n3884, A => n2024, ZN => n2017);
   U2065 : OAI22_X1 port map( A1 => n553, A2 => n1855, B1 => n521, B2 => n1856,
                           ZN => n2024);
   U2066 : NAND4_X1 port map( A1 => n2025, A2 => n2026, A3 => n2027, A4 => 
                           n2028, ZN => n2015);
   U2067 : AOI221_X1 port map( B1 => n1861, B2 => n3916, C1 => n1862, C2 => 
                           n3948, A => n2029, ZN => n2028);
   U2068 : OAI22_X1 port map( A1 => n425, A2 => n1864, B1 => n393, B2 => n1865,
                           ZN => n2029);
   U2069 : AOI221_X1 port map( B1 => n1866, B2 => n3980, C1 => n1867, C2 => 
                           n4012, A => n2030, ZN => n2027);
   U2070 : OAI22_X1 port map( A1 => n297, A2 => n1869, B1 => n265, B2 => n1870,
                           ZN => n2030);
   U2071 : AOI221_X1 port map( B1 => n1871, B2 => n145, C1 => n1872, C2 => n17,
                           A => n2031, ZN => n2026);
   U2072 : OAI22_X1 port map( A1 => n81, A2 => n1874, B1 => n209, B2 => n1875, 
                           ZN => n2031);
   U2073 : AOI221_X1 port map( B1 => n1876, B2 => n146, C1 => n1877, C2 => n18,
                           A => n2032, ZN => n2025);
   U2074 : OAI22_X1 port map( A1 => n82, A2 => n1879, B1 => n210, B2 => n1880, 
                           ZN => n2032);
   U2075 : OAI22_X1 port map( A1 => n2507, A2 => n1828, B1 => n2033, B2 => 
                           n1830, ZN => n2549);
   U2076 : NOR2_X1 port map( A1 => n2034, A2 => n2035, ZN => n2033);
   U2077 : NAND4_X1 port map( A1 => n2036, A2 => n2037, A3 => n2038, A4 => 
                           n2039, ZN => n2035);
   U2078 : AOI221_X1 port map( B1 => n1837, B2 => n3659, C1 => n1838, C2 => 
                           n3691, A => n2040, ZN => n2039);
   U2079 : OAI22_X1 port map( A1 => n1002, A2 => n1840, B1 => n970, B2 => n1841
                           , ZN => n2040);
   U2080 : AOI221_X1 port map( B1 => n1842, B2 => n3723, C1 => n1843, C2 => 
                           n3755, A => n2041, ZN => n2038);
   U2081 : OAI22_X1 port map( A1 => n874, A2 => n1845, B1 => n842, B2 => n1846,
                           ZN => n2041);
   U2082 : AOI221_X1 port map( B1 => n1847, B2 => n3787, C1 => n1848, C2 => 
                           n3819, A => n2042, ZN => n2037);
   U2083 : OAI22_X1 port map( A1 => n682, A2 => n1850, B1 => n650, B2 => n1851,
                           ZN => n2042);
   U2084 : AOI221_X1 port map( B1 => n1852, B2 => n3851, C1 => n1853, C2 => 
                           n3883, A => n2043, ZN => n2036);
   U2085 : OAI22_X1 port map( A1 => n554, A2 => n1855, B1 => n522, B2 => n1856,
                           ZN => n2043);
   U2086 : NAND4_X1 port map( A1 => n2044, A2 => n2045, A3 => n2046, A4 => 
                           n2047, ZN => n2034);
   U2087 : AOI221_X1 port map( B1 => n1861, B2 => n3915, C1 => n1862, C2 => 
                           n3947, A => n2048, ZN => n2047);
   U2088 : OAI22_X1 port map( A1 => n426, A2 => n1864, B1 => n394, B2 => n1865,
                           ZN => n2048);
   U2089 : AOI221_X1 port map( B1 => n1866, B2 => n3979, C1 => n1867, C2 => 
                           n4011, A => n2049, ZN => n2046);
   U2090 : OAI22_X1 port map( A1 => n298, A2 => n1869, B1 => n266, B2 => n1870,
                           ZN => n2049);
   U2091 : AOI221_X1 port map( B1 => n1871, B2 => n147, C1 => n1872, C2 => n19,
                           A => n2050, ZN => n2045);
   U2092 : OAI22_X1 port map( A1 => n83, A2 => n1874, B1 => n211, B2 => n1875, 
                           ZN => n2050);
   U2093 : AOI221_X1 port map( B1 => n1876, B2 => n148, C1 => n1877, C2 => n20,
                           A => n2051, ZN => n2044);
   U2094 : OAI22_X1 port map( A1 => n84, A2 => n1879, B1 => n212, B2 => n1880, 
                           ZN => n2051);
   U2095 : OAI22_X1 port map( A1 => n2506, A2 => n1828, B1 => n2052, B2 => 
                           n1830, ZN => n2548);
   U2096 : NOR2_X1 port map( A1 => n2053, A2 => n2054, ZN => n2052);
   U2097 : NAND4_X1 port map( A1 => n2055, A2 => n2056, A3 => n2057, A4 => 
                           n2058, ZN => n2054);
   U2098 : AOI221_X1 port map( B1 => n1837, B2 => n3658, C1 => n1838, C2 => 
                           n3690, A => n2059, ZN => n2058);
   U2099 : OAI22_X1 port map( A1 => n1003, A2 => n1840, B1 => n971, B2 => n1841
                           , ZN => n2059);
   U2100 : AOI221_X1 port map( B1 => n1842, B2 => n3722, C1 => n1843, C2 => 
                           n3754, A => n2060, ZN => n2057);
   U2101 : OAI22_X1 port map( A1 => n875, A2 => n1845, B1 => n843, B2 => n1846,
                           ZN => n2060);
   U2102 : AOI221_X1 port map( B1 => n1847, B2 => n3786, C1 => n1848, C2 => 
                           n3818, A => n2061, ZN => n2056);
   U2103 : OAI22_X1 port map( A1 => n683, A2 => n1850, B1 => n651, B2 => n1851,
                           ZN => n2061);
   U2104 : AOI221_X1 port map( B1 => n1852, B2 => n3850, C1 => n1853, C2 => 
                           n3882, A => n2062, ZN => n2055);
   U2105 : OAI22_X1 port map( A1 => n555, A2 => n1855, B1 => n523, B2 => n1856,
                           ZN => n2062);
   U2106 : NAND4_X1 port map( A1 => n2063, A2 => n2064, A3 => n2065, A4 => 
                           n2066, ZN => n2053);
   U2107 : AOI221_X1 port map( B1 => n1861, B2 => n3914, C1 => n1862, C2 => 
                           n3946, A => n2067, ZN => n2066);
   U2108 : OAI22_X1 port map( A1 => n427, A2 => n1864, B1 => n395, B2 => n1865,
                           ZN => n2067);
   U2109 : AOI221_X1 port map( B1 => n1866, B2 => n3978, C1 => n1867, C2 => 
                           n4010, A => n2068, ZN => n2065);
   U2110 : OAI22_X1 port map( A1 => n299, A2 => n1869, B1 => n267, B2 => n1870,
                           ZN => n2068);
   U2111 : AOI221_X1 port map( B1 => n1871, B2 => n149, C1 => n1872, C2 => n21,
                           A => n2069, ZN => n2064);
   U2112 : OAI22_X1 port map( A1 => n85, A2 => n1874, B1 => n213, B2 => n1875, 
                           ZN => n2069);
   U2113 : AOI221_X1 port map( B1 => n1876, B2 => n150, C1 => n1877, C2 => n22,
                           A => n2070, ZN => n2063);
   U2114 : OAI22_X1 port map( A1 => n86, A2 => n1879, B1 => n214, B2 => n1880, 
                           ZN => n2070);
   U2115 : OAI22_X1 port map( A1 => n2505, A2 => n1828, B1 => n2071, B2 => 
                           n1830, ZN => n2547);
   U2116 : NOR2_X1 port map( A1 => n2072, A2 => n2073, ZN => n2071);
   U2117 : NAND4_X1 port map( A1 => n2074, A2 => n2075, A3 => n2076, A4 => 
                           n2077, ZN => n2073);
   U2118 : AOI221_X1 port map( B1 => n1837, B2 => n3657, C1 => n1838, C2 => 
                           n3689, A => n2078, ZN => n2077);
   U2119 : OAI22_X1 port map( A1 => n1004, A2 => n1840, B1 => n972, B2 => n1841
                           , ZN => n2078);
   U2120 : AOI221_X1 port map( B1 => n1842, B2 => n3721, C1 => n1843, C2 => 
                           n3753, A => n2079, ZN => n2076);
   U2121 : OAI22_X1 port map( A1 => n876, A2 => n1845, B1 => n844, B2 => n1846,
                           ZN => n2079);
   U2122 : AOI221_X1 port map( B1 => n1847, B2 => n3785, C1 => n1848, C2 => 
                           n3817, A => n2080, ZN => n2075);
   U2123 : OAI22_X1 port map( A1 => n684, A2 => n1850, B1 => n652, B2 => n1851,
                           ZN => n2080);
   U2124 : AOI221_X1 port map( B1 => n1852, B2 => n3849, C1 => n1853, C2 => 
                           n3881, A => n2081, ZN => n2074);
   U2125 : OAI22_X1 port map( A1 => n556, A2 => n1855, B1 => n524, B2 => n1856,
                           ZN => n2081);
   U2126 : NAND4_X1 port map( A1 => n2082, A2 => n2083, A3 => n2084, A4 => 
                           n2085, ZN => n2072);
   U2127 : AOI221_X1 port map( B1 => n1861, B2 => n3913, C1 => n1862, C2 => 
                           n3945, A => n2086, ZN => n2085);
   U2128 : OAI22_X1 port map( A1 => n428, A2 => n1864, B1 => n396, B2 => n1865,
                           ZN => n2086);
   U2129 : AOI221_X1 port map( B1 => n1866, B2 => n3977, C1 => n1867, C2 => 
                           n4009, A => n2087, ZN => n2084);
   U2130 : OAI22_X1 port map( A1 => n300, A2 => n1869, B1 => n268, B2 => n1870,
                           ZN => n2087);
   U2131 : AOI221_X1 port map( B1 => n1871, B2 => n151, C1 => n1872, C2 => n23,
                           A => n2088, ZN => n2083);
   U2132 : OAI22_X1 port map( A1 => n87, A2 => n1874, B1 => n215, B2 => n1875, 
                           ZN => n2088);
   U2133 : AOI221_X1 port map( B1 => n1876, B2 => n152, C1 => n1877, C2 => n24,
                           A => n2089, ZN => n2082);
   U2134 : OAI22_X1 port map( A1 => n88, A2 => n1879, B1 => n216, B2 => n1880, 
                           ZN => n2089);
   U2135 : OAI22_X1 port map( A1 => n2504, A2 => n1828, B1 => n2090, B2 => 
                           n1830, ZN => n2546);
   U2136 : NOR2_X1 port map( A1 => n2091, A2 => n2092, ZN => n2090);
   U2137 : NAND4_X1 port map( A1 => n2093, A2 => n2094, A3 => n2095, A4 => 
                           n2096, ZN => n2092);
   U2138 : AOI221_X1 port map( B1 => n1837, B2 => n3656, C1 => n1838, C2 => 
                           n3688, A => n2097, ZN => n2096);
   U2139 : OAI22_X1 port map( A1 => n1005, A2 => n1840, B1 => n973, B2 => n1841
                           , ZN => n2097);
   U2140 : AOI221_X1 port map( B1 => n1842, B2 => n3720, C1 => n1843, C2 => 
                           n3752, A => n2098, ZN => n2095);
   U2141 : OAI22_X1 port map( A1 => n877, A2 => n1845, B1 => n845, B2 => n1846,
                           ZN => n2098);
   U2142 : AOI221_X1 port map( B1 => n1847, B2 => n3784, C1 => n1848, C2 => 
                           n3816, A => n2099, ZN => n2094);
   U2143 : OAI22_X1 port map( A1 => n685, A2 => n1850, B1 => n653, B2 => n1851,
                           ZN => n2099);
   U2144 : AOI221_X1 port map( B1 => n1852, B2 => n3848, C1 => n1853, C2 => 
                           n3880, A => n2100, ZN => n2093);
   U2145 : OAI22_X1 port map( A1 => n557, A2 => n1855, B1 => n525, B2 => n1856,
                           ZN => n2100);
   U2146 : NAND4_X1 port map( A1 => n2101, A2 => n2102, A3 => n2103, A4 => 
                           n2104, ZN => n2091);
   U2147 : AOI221_X1 port map( B1 => n1861, B2 => n3912, C1 => n1862, C2 => 
                           n3944, A => n2105, ZN => n2104);
   U2148 : OAI22_X1 port map( A1 => n429, A2 => n1864, B1 => n397, B2 => n1865,
                           ZN => n2105);
   U2149 : AOI221_X1 port map( B1 => n1866, B2 => n3976, C1 => n1867, C2 => 
                           n4008, A => n2106, ZN => n2103);
   U2150 : OAI22_X1 port map( A1 => n301, A2 => n1869, B1 => n269, B2 => n1870,
                           ZN => n2106);
   U2151 : AOI221_X1 port map( B1 => n1871, B2 => n153, C1 => n1872, C2 => n25,
                           A => n2107, ZN => n2102);
   U2152 : OAI22_X1 port map( A1 => n89, A2 => n1874, B1 => n217, B2 => n1875, 
                           ZN => n2107);
   U2153 : AOI221_X1 port map( B1 => n1876, B2 => n154, C1 => n1877, C2 => n26,
                           A => n2108, ZN => n2101);
   U2154 : OAI22_X1 port map( A1 => n90, A2 => n1879, B1 => n218, B2 => n1880, 
                           ZN => n2108);
   U2155 : OAI22_X1 port map( A1 => n2503, A2 => n1828, B1 => n2109, B2 => 
                           n1830, ZN => n2545);
   U2156 : NOR2_X1 port map( A1 => n2110, A2 => n2111, ZN => n2109);
   U2157 : NAND4_X1 port map( A1 => n2112, A2 => n2113, A3 => n2114, A4 => 
                           n2115, ZN => n2111);
   U2158 : AOI221_X1 port map( B1 => n1837, B2 => n3655, C1 => n1838, C2 => 
                           n3687, A => n2116, ZN => n2115);
   U2159 : OAI22_X1 port map( A1 => n1006, A2 => n1840, B1 => n974, B2 => n1841
                           , ZN => n2116);
   U2160 : AOI221_X1 port map( B1 => n1842, B2 => n3719, C1 => n1843, C2 => 
                           n3751, A => n2117, ZN => n2114);
   U2161 : OAI22_X1 port map( A1 => n878, A2 => n1845, B1 => n846, B2 => n1846,
                           ZN => n2117);
   U2162 : AOI221_X1 port map( B1 => n1847, B2 => n3783, C1 => n1848, C2 => 
                           n3815, A => n2118, ZN => n2113);
   U2163 : OAI22_X1 port map( A1 => n686, A2 => n1850, B1 => n654, B2 => n1851,
                           ZN => n2118);
   U2164 : AOI221_X1 port map( B1 => n1852, B2 => n3847, C1 => n1853, C2 => 
                           n3879, A => n2119, ZN => n2112);
   U2165 : OAI22_X1 port map( A1 => n558, A2 => n1855, B1 => n526, B2 => n1856,
                           ZN => n2119);
   U2166 : NAND4_X1 port map( A1 => n2120, A2 => n2121, A3 => n2122, A4 => 
                           n2123, ZN => n2110);
   U2167 : AOI221_X1 port map( B1 => n1861, B2 => n3911, C1 => n1862, C2 => 
                           n3943, A => n2124, ZN => n2123);
   U2168 : OAI22_X1 port map( A1 => n430, A2 => n1864, B1 => n398, B2 => n1865,
                           ZN => n2124);
   U2169 : AOI221_X1 port map( B1 => n1866, B2 => n3975, C1 => n1867, C2 => 
                           n4007, A => n2125, ZN => n2122);
   U2170 : OAI22_X1 port map( A1 => n302, A2 => n1869, B1 => n270, B2 => n1870,
                           ZN => n2125);
   U2171 : AOI221_X1 port map( B1 => n1871, B2 => n155, C1 => n1872, C2 => n27,
                           A => n2126, ZN => n2121);
   U2172 : OAI22_X1 port map( A1 => n91, A2 => n1874, B1 => n219, B2 => n1875, 
                           ZN => n2126);
   U2173 : AOI221_X1 port map( B1 => n1876, B2 => n156, C1 => n1877, C2 => n28,
                           A => n2127, ZN => n2120);
   U2174 : OAI22_X1 port map( A1 => n92, A2 => n1879, B1 => n220, B2 => n1880, 
                           ZN => n2127);
   U2175 : OAI22_X1 port map( A1 => n2502, A2 => n1828, B1 => n2128, B2 => 
                           n1830, ZN => n2544);
   U2176 : NOR2_X1 port map( A1 => n2129, A2 => n2130, ZN => n2128);
   U2177 : NAND4_X1 port map( A1 => n2131, A2 => n2132, A3 => n2133, A4 => 
                           n2134, ZN => n2130);
   U2178 : AOI221_X1 port map( B1 => n1837, B2 => n3654, C1 => n1838, C2 => 
                           n3686, A => n2135, ZN => n2134);
   U2179 : OAI22_X1 port map( A1 => n1007, A2 => n1840, B1 => n975, B2 => n1841
                           , ZN => n2135);
   U2180 : AOI221_X1 port map( B1 => n1842, B2 => n3718, C1 => n1843, C2 => 
                           n3750, A => n2136, ZN => n2133);
   U2181 : OAI22_X1 port map( A1 => n879, A2 => n1845, B1 => n847, B2 => n1846,
                           ZN => n2136);
   U2182 : AOI221_X1 port map( B1 => n1847, B2 => n3782, C1 => n1848, C2 => 
                           n3814, A => n2137, ZN => n2132);
   U2183 : OAI22_X1 port map( A1 => n687, A2 => n1850, B1 => n655, B2 => n1851,
                           ZN => n2137);
   U2184 : AOI221_X1 port map( B1 => n1852, B2 => n3846, C1 => n1853, C2 => 
                           n3878, A => n2138, ZN => n2131);
   U2185 : OAI22_X1 port map( A1 => n559, A2 => n1855, B1 => n527, B2 => n1856,
                           ZN => n2138);
   U2186 : NAND4_X1 port map( A1 => n2139, A2 => n2140, A3 => n2141, A4 => 
                           n2142, ZN => n2129);
   U2187 : AOI221_X1 port map( B1 => n1861, B2 => n3910, C1 => n1862, C2 => 
                           n3942, A => n2143, ZN => n2142);
   U2188 : OAI22_X1 port map( A1 => n431, A2 => n1864, B1 => n399, B2 => n1865,
                           ZN => n2143);
   U2189 : AOI221_X1 port map( B1 => n1866, B2 => n3974, C1 => n1867, C2 => 
                           n4006, A => n2144, ZN => n2141);
   U2190 : OAI22_X1 port map( A1 => n303, A2 => n1869, B1 => n271, B2 => n1870,
                           ZN => n2144);
   U2191 : AOI221_X1 port map( B1 => n1871, B2 => n157, C1 => n1872, C2 => n29,
                           A => n2145, ZN => n2140);
   U2192 : OAI22_X1 port map( A1 => n93, A2 => n1874, B1 => n221, B2 => n1875, 
                           ZN => n2145);
   U2193 : AOI221_X1 port map( B1 => n1876, B2 => n158, C1 => n1877, C2 => n30,
                           A => n2146, ZN => n2139);
   U2194 : OAI22_X1 port map( A1 => n94, A2 => n1879, B1 => n222, B2 => n1880, 
                           ZN => n2146);
   U2195 : OAI22_X1 port map( A1 => n2501, A2 => n1828, B1 => n2147, B2 => 
                           n1830, ZN => n2543);
   U2196 : NOR2_X1 port map( A1 => n2148, A2 => n2149, ZN => n2147);
   U2197 : NAND4_X1 port map( A1 => n2150, A2 => n2151, A3 => n2152, A4 => 
                           n2153, ZN => n2149);
   U2198 : AOI221_X1 port map( B1 => n1837, B2 => n3653, C1 => n1838, C2 => 
                           n3685, A => n2154, ZN => n2153);
   U2199 : OAI22_X1 port map( A1 => n1008, A2 => n1840, B1 => n976, B2 => n1841
                           , ZN => n2154);
   U2200 : AOI221_X1 port map( B1 => n1842, B2 => n3717, C1 => n1843, C2 => 
                           n3749, A => n2155, ZN => n2152);
   U2201 : OAI22_X1 port map( A1 => n880, A2 => n1845, B1 => n848, B2 => n1846,
                           ZN => n2155);
   U2202 : AOI221_X1 port map( B1 => n1847, B2 => n3781, C1 => n1848, C2 => 
                           n3813, A => n2156, ZN => n2151);
   U2203 : OAI22_X1 port map( A1 => n688, A2 => n1850, B1 => n656, B2 => n1851,
                           ZN => n2156);
   U2204 : AOI221_X1 port map( B1 => n1852, B2 => n3845, C1 => n1853, C2 => 
                           n3877, A => n2157, ZN => n2150);
   U2205 : OAI22_X1 port map( A1 => n560, A2 => n1855, B1 => n528, B2 => n1856,
                           ZN => n2157);
   U2206 : NAND4_X1 port map( A1 => n2158, A2 => n2159, A3 => n2160, A4 => 
                           n2161, ZN => n2148);
   U2207 : AOI221_X1 port map( B1 => n1861, B2 => n3909, C1 => n1862, C2 => 
                           n3941, A => n2162, ZN => n2161);
   U2208 : OAI22_X1 port map( A1 => n432, A2 => n1864, B1 => n400, B2 => n1865,
                           ZN => n2162);
   U2209 : AOI221_X1 port map( B1 => n1866, B2 => n3973, C1 => n1867, C2 => 
                           n4005, A => n2163, ZN => n2160);
   U2210 : OAI22_X1 port map( A1 => n304, A2 => n1869, B1 => n272, B2 => n1870,
                           ZN => n2163);
   U2211 : AOI221_X1 port map( B1 => n1871, B2 => n159, C1 => n1872, C2 => n31,
                           A => n2164, ZN => n2159);
   U2212 : OAI22_X1 port map( A1 => n95, A2 => n1874, B1 => n223, B2 => n1875, 
                           ZN => n2164);
   U2213 : AOI221_X1 port map( B1 => n1876, B2 => n160, C1 => n1877, C2 => n32,
                           A => n2165, ZN => n2158);
   U2214 : OAI22_X1 port map( A1 => n96, A2 => n1879, B1 => n224, B2 => n1880, 
                           ZN => n2165);
   U2215 : OAI22_X1 port map( A1 => n2500, A2 => n1828, B1 => n2166, B2 => 
                           n1830, ZN => n2542);
   U2216 : NOR2_X1 port map( A1 => n2167, A2 => n2168, ZN => n2166);
   U2217 : NAND4_X1 port map( A1 => n2169, A2 => n2170, A3 => n2171, A4 => 
                           n2172, ZN => n2168);
   U2218 : AOI221_X1 port map( B1 => n1837, B2 => n3652, C1 => n1838, C2 => 
                           n3684, A => n2173, ZN => n2172);
   U2219 : OAI22_X1 port map( A1 => n1009, A2 => n1840, B1 => n977, B2 => n1841
                           , ZN => n2173);
   U2220 : AOI221_X1 port map( B1 => n1842, B2 => n3716, C1 => n1843, C2 => 
                           n3748, A => n2174, ZN => n2171);
   U2221 : OAI22_X1 port map( A1 => n881, A2 => n1845, B1 => n849, B2 => n1846,
                           ZN => n2174);
   U2222 : AOI221_X1 port map( B1 => n1847, B2 => n3780, C1 => n1848, C2 => 
                           n3812, A => n2175, ZN => n2170);
   U2223 : OAI22_X1 port map( A1 => n689, A2 => n1850, B1 => n657, B2 => n1851,
                           ZN => n2175);
   U2224 : AOI221_X1 port map( B1 => n1852, B2 => n3844, C1 => n1853, C2 => 
                           n3876, A => n2176, ZN => n2169);
   U2225 : OAI22_X1 port map( A1 => n561, A2 => n1855, B1 => n529, B2 => n1856,
                           ZN => n2176);
   U2226 : NAND4_X1 port map( A1 => n2177, A2 => n2178, A3 => n2179, A4 => 
                           n2180, ZN => n2167);
   U2227 : AOI221_X1 port map( B1 => n1861, B2 => n3908, C1 => n1862, C2 => 
                           n3940, A => n2181, ZN => n2180);
   U2228 : OAI22_X1 port map( A1 => n433, A2 => n1864, B1 => n401, B2 => n1865,
                           ZN => n2181);
   U2229 : AOI221_X1 port map( B1 => n1866, B2 => n3972, C1 => n1867, C2 => 
                           n4004, A => n2182, ZN => n2179);
   U2230 : OAI22_X1 port map( A1 => n305, A2 => n1869, B1 => n273, B2 => n1870,
                           ZN => n2182);
   U2231 : AOI221_X1 port map( B1 => n1871, B2 => n161, C1 => n1872, C2 => n33,
                           A => n2183, ZN => n2178);
   U2232 : OAI22_X1 port map( A1 => n97, A2 => n1874, B1 => n225, B2 => n1875, 
                           ZN => n2183);
   U2233 : AOI221_X1 port map( B1 => n1876, B2 => n162, C1 => n1877, C2 => n34,
                           A => n2184, ZN => n2177);
   U2234 : OAI22_X1 port map( A1 => n98, A2 => n1879, B1 => n226, B2 => n1880, 
                           ZN => n2184);
   U2235 : OAI22_X1 port map( A1 => n2499, A2 => n1828, B1 => n2185, B2 => 
                           n1830, ZN => n2541);
   U2236 : NOR2_X1 port map( A1 => n2186, A2 => n2187, ZN => n2185);
   U2237 : NAND4_X1 port map( A1 => n2188, A2 => n2189, A3 => n2190, A4 => 
                           n2191, ZN => n2187);
   U2238 : AOI221_X1 port map( B1 => n1837, B2 => n3651, C1 => n1838, C2 => 
                           n3683, A => n2192, ZN => n2191);
   U2239 : OAI22_X1 port map( A1 => n1010, A2 => n1840, B1 => n978, B2 => n1841
                           , ZN => n2192);
   U2240 : AOI221_X1 port map( B1 => n1842, B2 => n3715, C1 => n1843, C2 => 
                           n3747, A => n2193, ZN => n2190);
   U2241 : OAI22_X1 port map( A1 => n882, A2 => n1845, B1 => n850, B2 => n1846,
                           ZN => n2193);
   U2242 : AOI221_X1 port map( B1 => n1847, B2 => n3779, C1 => n1848, C2 => 
                           n3811, A => n2194, ZN => n2189);
   U2243 : OAI22_X1 port map( A1 => n690, A2 => n1850, B1 => n658, B2 => n1851,
                           ZN => n2194);
   U2244 : AOI221_X1 port map( B1 => n1852, B2 => n3843, C1 => n1853, C2 => 
                           n3875, A => n2195, ZN => n2188);
   U2245 : OAI22_X1 port map( A1 => n562, A2 => n1855, B1 => n530, B2 => n1856,
                           ZN => n2195);
   U2246 : NAND4_X1 port map( A1 => n2196, A2 => n2197, A3 => n2198, A4 => 
                           n2199, ZN => n2186);
   U2247 : AOI221_X1 port map( B1 => n1861, B2 => n3907, C1 => n1862, C2 => 
                           n3939, A => n2200, ZN => n2199);
   U2248 : OAI22_X1 port map( A1 => n434, A2 => n1864, B1 => n402, B2 => n1865,
                           ZN => n2200);
   U2249 : AOI221_X1 port map( B1 => n1866, B2 => n3971, C1 => n1867, C2 => 
                           n4003, A => n2201, ZN => n2198);
   U2250 : OAI22_X1 port map( A1 => n306, A2 => n1869, B1 => n274, B2 => n1870,
                           ZN => n2201);
   U2251 : AOI221_X1 port map( B1 => n1871, B2 => n163, C1 => n1872, C2 => n35,
                           A => n2202, ZN => n2197);
   U2252 : OAI22_X1 port map( A1 => n99, A2 => n1874, B1 => n227, B2 => n1875, 
                           ZN => n2202);
   U2253 : AOI221_X1 port map( B1 => n1876, B2 => n164, C1 => n1877, C2 => n36,
                           A => n2203, ZN => n2196);
   U2254 : OAI22_X1 port map( A1 => n100, A2 => n1879, B1 => n228, B2 => n1880,
                           ZN => n2203);
   U2255 : OAI22_X1 port map( A1 => n2498, A2 => n1828, B1 => n2204, B2 => 
                           n1830, ZN => n2540);
   U2256 : NOR2_X1 port map( A1 => n2205, A2 => n2206, ZN => n2204);
   U2257 : NAND4_X1 port map( A1 => n2207, A2 => n2208, A3 => n2209, A4 => 
                           n2210, ZN => n2206);
   U2258 : AOI221_X1 port map( B1 => n1837, B2 => n3650, C1 => n1838, C2 => 
                           n3682, A => n2211, ZN => n2210);
   U2259 : OAI22_X1 port map( A1 => n1011, A2 => n1840, B1 => n979, B2 => n1841
                           , ZN => n2211);
   U2260 : AOI221_X1 port map( B1 => n1842, B2 => n3714, C1 => n1843, C2 => 
                           n3746, A => n2212, ZN => n2209);
   U2261 : OAI22_X1 port map( A1 => n883, A2 => n1845, B1 => n851, B2 => n1846,
                           ZN => n2212);
   U2262 : AOI221_X1 port map( B1 => n1847, B2 => n3778, C1 => n1848, C2 => 
                           n3810, A => n2213, ZN => n2208);
   U2263 : OAI22_X1 port map( A1 => n691, A2 => n1850, B1 => n659, B2 => n1851,
                           ZN => n2213);
   U2264 : AOI221_X1 port map( B1 => n1852, B2 => n3842, C1 => n1853, C2 => 
                           n3874, A => n2214, ZN => n2207);
   U2265 : OAI22_X1 port map( A1 => n563, A2 => n1855, B1 => n531, B2 => n1856,
                           ZN => n2214);
   U2266 : NAND4_X1 port map( A1 => n2215, A2 => n2216, A3 => n2217, A4 => 
                           n2218, ZN => n2205);
   U2267 : AOI221_X1 port map( B1 => n1861, B2 => n3906, C1 => n1862, C2 => 
                           n3938, A => n2219, ZN => n2218);
   U2268 : OAI22_X1 port map( A1 => n435, A2 => n1864, B1 => n403, B2 => n1865,
                           ZN => n2219);
   U2269 : AOI221_X1 port map( B1 => n1866, B2 => n3970, C1 => n1867, C2 => 
                           n4002, A => n2220, ZN => n2217);
   U2270 : OAI22_X1 port map( A1 => n307, A2 => n1869, B1 => n275, B2 => n1870,
                           ZN => n2220);
   U2271 : AOI221_X1 port map( B1 => n1871, B2 => n165, C1 => n1872, C2 => n37,
                           A => n2221, ZN => n2216);
   U2272 : OAI22_X1 port map( A1 => n101, A2 => n1874, B1 => n229, B2 => n1875,
                           ZN => n2221);
   U2273 : AOI221_X1 port map( B1 => n1876, B2 => n166, C1 => n1877, C2 => n38,
                           A => n2222, ZN => n2215);
   U2274 : OAI22_X1 port map( A1 => n102, A2 => n1879, B1 => n230, B2 => n1880,
                           ZN => n2222);
   U2275 : OAI22_X1 port map( A1 => n2497, A2 => n1828, B1 => n2223, B2 => 
                           n1830, ZN => n2539);
   U2276 : NOR2_X1 port map( A1 => n2224, A2 => n2225, ZN => n2223);
   U2277 : NAND4_X1 port map( A1 => n2226, A2 => n2227, A3 => n2228, A4 => 
                           n2229, ZN => n2225);
   U2278 : AOI221_X1 port map( B1 => n1837, B2 => n3649, C1 => n1838, C2 => 
                           n3681, A => n2230, ZN => n2229);
   U2279 : OAI22_X1 port map( A1 => n1012, A2 => n1840, B1 => n980, B2 => n1841
                           , ZN => n2230);
   U2280 : AOI221_X1 port map( B1 => n1842, B2 => n3713, C1 => n1843, C2 => 
                           n3745, A => n2231, ZN => n2228);
   U2281 : OAI22_X1 port map( A1 => n884, A2 => n1845, B1 => n852, B2 => n1846,
                           ZN => n2231);
   U2282 : AOI221_X1 port map( B1 => n1847, B2 => n3777, C1 => n1848, C2 => 
                           n3809, A => n2232, ZN => n2227);
   U2283 : OAI22_X1 port map( A1 => n692, A2 => n1850, B1 => n660, B2 => n1851,
                           ZN => n2232);
   U2284 : AOI221_X1 port map( B1 => n1852, B2 => n3841, C1 => n1853, C2 => 
                           n3873, A => n2233, ZN => n2226);
   U2285 : OAI22_X1 port map( A1 => n564, A2 => n1855, B1 => n532, B2 => n1856,
                           ZN => n2233);
   U2286 : NAND4_X1 port map( A1 => n2234, A2 => n2235, A3 => n2236, A4 => 
                           n2237, ZN => n2224);
   U2287 : AOI221_X1 port map( B1 => n1861, B2 => n3905, C1 => n1862, C2 => 
                           n3937, A => n2238, ZN => n2237);
   U2288 : OAI22_X1 port map( A1 => n436, A2 => n1864, B1 => n404, B2 => n1865,
                           ZN => n2238);
   U2289 : AOI221_X1 port map( B1 => n1866, B2 => n3969, C1 => n1867, C2 => 
                           n4001, A => n2239, ZN => n2236);
   U2290 : OAI22_X1 port map( A1 => n308, A2 => n1869, B1 => n276, B2 => n1870,
                           ZN => n2239);
   U2291 : AOI221_X1 port map( B1 => n1871, B2 => n167, C1 => n1872, C2 => n39,
                           A => n2240, ZN => n2235);
   U2292 : OAI22_X1 port map( A1 => n103, A2 => n1874, B1 => n231, B2 => n1875,
                           ZN => n2240);
   U2293 : AOI221_X1 port map( B1 => n1876, B2 => n168, C1 => n1877, C2 => n40,
                           A => n2241, ZN => n2234);
   U2294 : OAI22_X1 port map( A1 => n104, A2 => n1879, B1 => n232, B2 => n1880,
                           ZN => n2241);
   U2295 : OAI22_X1 port map( A1 => n2496, A2 => n1828, B1 => n2242, B2 => 
                           n1830, ZN => n2538);
   U2296 : NOR2_X1 port map( A1 => n2243, A2 => n2244, ZN => n2242);
   U2297 : NAND4_X1 port map( A1 => n2245, A2 => n2246, A3 => n2247, A4 => 
                           n2248, ZN => n2244);
   U2298 : AOI221_X1 port map( B1 => n1837, B2 => n3648, C1 => n1838, C2 => 
                           n3680, A => n2249, ZN => n2248);
   U2299 : OAI22_X1 port map( A1 => n1013, A2 => n1840, B1 => n981, B2 => n1841
                           , ZN => n2249);
   U2300 : AOI221_X1 port map( B1 => n1842, B2 => n3712, C1 => n1843, C2 => 
                           n3744, A => n2250, ZN => n2247);
   U2301 : OAI22_X1 port map( A1 => n885, A2 => n1845, B1 => n853, B2 => n1846,
                           ZN => n2250);
   U2302 : AOI221_X1 port map( B1 => n1847, B2 => n3776, C1 => n1848, C2 => 
                           n3808, A => n2251, ZN => n2246);
   U2303 : OAI22_X1 port map( A1 => n693, A2 => n1850, B1 => n661, B2 => n1851,
                           ZN => n2251);
   U2304 : AOI221_X1 port map( B1 => n1852, B2 => n3840, C1 => n1853, C2 => 
                           n3872, A => n2252, ZN => n2245);
   U2305 : OAI22_X1 port map( A1 => n565, A2 => n1855, B1 => n533, B2 => n1856,
                           ZN => n2252);
   U2306 : NAND4_X1 port map( A1 => n2253, A2 => n2254, A3 => n2255, A4 => 
                           n2256, ZN => n2243);
   U2307 : AOI221_X1 port map( B1 => n1861, B2 => n3904, C1 => n1862, C2 => 
                           n3936, A => n2257, ZN => n2256);
   U2308 : OAI22_X1 port map( A1 => n437, A2 => n1864, B1 => n405, B2 => n1865,
                           ZN => n2257);
   U2309 : AOI221_X1 port map( B1 => n1866, B2 => n3968, C1 => n1867, C2 => 
                           n4000, A => n2258, ZN => n2255);
   U2310 : OAI22_X1 port map( A1 => n309, A2 => n1869, B1 => n277, B2 => n1870,
                           ZN => n2258);
   U2311 : AOI221_X1 port map( B1 => n1871, B2 => n169, C1 => n1872, C2 => n41,
                           A => n2259, ZN => n2254);
   U2312 : OAI22_X1 port map( A1 => n105, A2 => n1874, B1 => n233, B2 => n1875,
                           ZN => n2259);
   U2313 : AOI221_X1 port map( B1 => n1876, B2 => n170, C1 => n1877, C2 => n42,
                           A => n2260, ZN => n2253);
   U2314 : OAI22_X1 port map( A1 => n106, A2 => n1879, B1 => n234, B2 => n1880,
                           ZN => n2260);
   U2315 : OAI22_X1 port map( A1 => n2495, A2 => n1828, B1 => n2261, B2 => 
                           n1830, ZN => n2537);
   U2316 : NOR2_X1 port map( A1 => n2262, A2 => n2263, ZN => n2261);
   U2317 : NAND4_X1 port map( A1 => n2264, A2 => n2265, A3 => n2266, A4 => 
                           n2267, ZN => n2263);
   U2318 : AOI221_X1 port map( B1 => n1837, B2 => n3647, C1 => n1838, C2 => 
                           n3679, A => n2268, ZN => n2267);
   U2319 : OAI22_X1 port map( A1 => n1014, A2 => n1840, B1 => n982, B2 => n1841
                           , ZN => n2268);
   U2320 : AOI221_X1 port map( B1 => n1842, B2 => n3711, C1 => n1843, C2 => 
                           n3743, A => n2269, ZN => n2266);
   U2321 : OAI22_X1 port map( A1 => n886, A2 => n1845, B1 => n854, B2 => n1846,
                           ZN => n2269);
   U2322 : AOI221_X1 port map( B1 => n1847, B2 => n3775, C1 => n1848, C2 => 
                           n3807, A => n2270, ZN => n2265);
   U2323 : OAI22_X1 port map( A1 => n694, A2 => n1850, B1 => n662, B2 => n1851,
                           ZN => n2270);
   U2324 : AOI221_X1 port map( B1 => n1852, B2 => n3839, C1 => n1853, C2 => 
                           n3871, A => n2271, ZN => n2264);
   U2325 : OAI22_X1 port map( A1 => n566, A2 => n1855, B1 => n534, B2 => n1856,
                           ZN => n2271);
   U2326 : NAND4_X1 port map( A1 => n2272, A2 => n2273, A3 => n2274, A4 => 
                           n2275, ZN => n2262);
   U2327 : AOI221_X1 port map( B1 => n1861, B2 => n3903, C1 => n1862, C2 => 
                           n3935, A => n2276, ZN => n2275);
   U2328 : OAI22_X1 port map( A1 => n438, A2 => n1864, B1 => n406, B2 => n1865,
                           ZN => n2276);
   U2329 : AOI221_X1 port map( B1 => n1866, B2 => n3967, C1 => n1867, C2 => 
                           n3999, A => n2277, ZN => n2274);
   U2330 : OAI22_X1 port map( A1 => n310, A2 => n1869, B1 => n278, B2 => n1870,
                           ZN => n2277);
   U2331 : AOI221_X1 port map( B1 => n1871, B2 => n171, C1 => n1872, C2 => n43,
                           A => n2278, ZN => n2273);
   U2332 : OAI22_X1 port map( A1 => n107, A2 => n1874, B1 => n235, B2 => n1875,
                           ZN => n2278);
   U2333 : AOI221_X1 port map( B1 => n1876, B2 => n172, C1 => n1877, C2 => n44,
                           A => n2279, ZN => n2272);
   U2334 : OAI22_X1 port map( A1 => n108, A2 => n1879, B1 => n236, B2 => n1880,
                           ZN => n2279);
   U2335 : OAI22_X1 port map( A1 => n2494, A2 => n1828, B1 => n2280, B2 => 
                           n1830, ZN => n2536);
   U2336 : NOR2_X1 port map( A1 => n2281, A2 => n2282, ZN => n2280);
   U2337 : NAND4_X1 port map( A1 => n2283, A2 => n2284, A3 => n2285, A4 => 
                           n2286, ZN => n2282);
   U2338 : AOI221_X1 port map( B1 => n1837, B2 => n3646, C1 => n1838, C2 => 
                           n3678, A => n2287, ZN => n2286);
   U2339 : OAI22_X1 port map( A1 => n1015, A2 => n1840, B1 => n983, B2 => n1841
                           , ZN => n2287);
   U2340 : AOI221_X1 port map( B1 => n1842, B2 => n3710, C1 => n1843, C2 => 
                           n3742, A => n2288, ZN => n2285);
   U2341 : OAI22_X1 port map( A1 => n887, A2 => n1845, B1 => n855, B2 => n1846,
                           ZN => n2288);
   U2342 : AOI221_X1 port map( B1 => n1847, B2 => n3774, C1 => n1848, C2 => 
                           n3806, A => n2289, ZN => n2284);
   U2343 : OAI22_X1 port map( A1 => n695, A2 => n1850, B1 => n663, B2 => n1851,
                           ZN => n2289);
   U2344 : AOI221_X1 port map( B1 => n1852, B2 => n3838, C1 => n1853, C2 => 
                           n3870, A => n2290, ZN => n2283);
   U2345 : OAI22_X1 port map( A1 => n567, A2 => n1855, B1 => n535, B2 => n1856,
                           ZN => n2290);
   U2346 : NAND4_X1 port map( A1 => n2291, A2 => n2292, A3 => n2293, A4 => 
                           n2294, ZN => n2281);
   U2347 : AOI221_X1 port map( B1 => n1861, B2 => n3902, C1 => n1862, C2 => 
                           n3934, A => n2295, ZN => n2294);
   U2348 : OAI22_X1 port map( A1 => n439, A2 => n1864, B1 => n407, B2 => n1865,
                           ZN => n2295);
   U2349 : AOI221_X1 port map( B1 => n1866, B2 => n3966, C1 => n1867, C2 => 
                           n3998, A => n2296, ZN => n2293);
   U2350 : OAI22_X1 port map( A1 => n311, A2 => n1869, B1 => n279, B2 => n1870,
                           ZN => n2296);
   U2351 : AOI221_X1 port map( B1 => n1871, B2 => n173, C1 => n1872, C2 => n45,
                           A => n2297, ZN => n2292);
   U2352 : OAI22_X1 port map( A1 => n109, A2 => n1874, B1 => n237, B2 => n1875,
                           ZN => n2297);
   U2353 : AOI221_X1 port map( B1 => n1876, B2 => n174, C1 => n1877, C2 => n46,
                           A => n2298, ZN => n2291);
   U2354 : OAI22_X1 port map( A1 => n110, A2 => n1879, B1 => n238, B2 => n1880,
                           ZN => n2298);
   U2355 : OAI22_X1 port map( A1 => n2493, A2 => n1828, B1 => n2299, B2 => 
                           n1830, ZN => n2535);
   U2356 : NOR2_X1 port map( A1 => n2300, A2 => n2301, ZN => n2299);
   U2357 : NAND4_X1 port map( A1 => n2302, A2 => n2303, A3 => n2304, A4 => 
                           n2305, ZN => n2301);
   U2358 : AOI221_X1 port map( B1 => n1837, B2 => n3645, C1 => n1838, C2 => 
                           n3677, A => n2306, ZN => n2305);
   U2359 : OAI22_X1 port map( A1 => n1016, A2 => n1840, B1 => n984, B2 => n1841
                           , ZN => n2306);
   U2360 : AOI221_X1 port map( B1 => n1842, B2 => n3709, C1 => n1843, C2 => 
                           n3741, A => n2307, ZN => n2304);
   U2361 : OAI22_X1 port map( A1 => n888, A2 => n1845, B1 => n856, B2 => n1846,
                           ZN => n2307);
   U2362 : AOI221_X1 port map( B1 => n1847, B2 => n3773, C1 => n1848, C2 => 
                           n3805, A => n2308, ZN => n2303);
   U2363 : OAI22_X1 port map( A1 => n696, A2 => n1850, B1 => n664, B2 => n1851,
                           ZN => n2308);
   U2364 : AOI221_X1 port map( B1 => n1852, B2 => n3837, C1 => n1853, C2 => 
                           n3869, A => n2309, ZN => n2302);
   U2365 : OAI22_X1 port map( A1 => n568, A2 => n1855, B1 => n536, B2 => n1856,
                           ZN => n2309);
   U2366 : NAND4_X1 port map( A1 => n2310, A2 => n2311, A3 => n2312, A4 => 
                           n2313, ZN => n2300);
   U2367 : AOI221_X1 port map( B1 => n1861, B2 => n3901, C1 => n1862, C2 => 
                           n3933, A => n2314, ZN => n2313);
   U2368 : OAI22_X1 port map( A1 => n440, A2 => n1864, B1 => n408, B2 => n1865,
                           ZN => n2314);
   U2369 : AOI221_X1 port map( B1 => n1866, B2 => n3965, C1 => n1867, C2 => 
                           n3997, A => n2315, ZN => n2312);
   U2370 : OAI22_X1 port map( A1 => n312, A2 => n1869, B1 => n280, B2 => n1870,
                           ZN => n2315);
   U2371 : AOI221_X1 port map( B1 => n1871, B2 => n175, C1 => n1872, C2 => n47,
                           A => n2316, ZN => n2311);
   U2372 : OAI22_X1 port map( A1 => n111, A2 => n1874, B1 => n239, B2 => n1875,
                           ZN => n2316);
   U2373 : AOI221_X1 port map( B1 => n1876, B2 => n176, C1 => n1877, C2 => n48,
                           A => n2317, ZN => n2310);
   U2374 : OAI22_X1 port map( A1 => n112, A2 => n1879, B1 => n240, B2 => n1880,
                           ZN => n2317);
   U2375 : OAI22_X1 port map( A1 => n2492, A2 => n1828, B1 => n2318, B2 => 
                           n1830, ZN => n2534);
   U2376 : NOR2_X1 port map( A1 => n2319, A2 => n2320, ZN => n2318);
   U2377 : NAND4_X1 port map( A1 => n2321, A2 => n2322, A3 => n2323, A4 => 
                           n2324, ZN => n2320);
   U2378 : AOI221_X1 port map( B1 => n1837, B2 => n3644, C1 => n1838, C2 => 
                           n3676, A => n2325, ZN => n2324);
   U2379 : OAI22_X1 port map( A1 => n1017, A2 => n1840, B1 => n985, B2 => n1841
                           , ZN => n2325);
   U2380 : AOI221_X1 port map( B1 => n1842, B2 => n3708, C1 => n1843, C2 => 
                           n3740, A => n2326, ZN => n2323);
   U2381 : OAI22_X1 port map( A1 => n889, A2 => n1845, B1 => n857, B2 => n1846,
                           ZN => n2326);
   U2382 : AOI221_X1 port map( B1 => n1847, B2 => n3772, C1 => n1848, C2 => 
                           n3804, A => n2327, ZN => n2322);
   U2383 : OAI22_X1 port map( A1 => n697, A2 => n1850, B1 => n665, B2 => n1851,
                           ZN => n2327);
   U2384 : AOI221_X1 port map( B1 => n1852, B2 => n3836, C1 => n1853, C2 => 
                           n3868, A => n2328, ZN => n2321);
   U2385 : OAI22_X1 port map( A1 => n569, A2 => n1855, B1 => n537, B2 => n1856,
                           ZN => n2328);
   U2386 : NAND4_X1 port map( A1 => n2329, A2 => n2330, A3 => n2331, A4 => 
                           n2332, ZN => n2319);
   U2387 : AOI221_X1 port map( B1 => n1861, B2 => n3900, C1 => n1862, C2 => 
                           n3932, A => n2333, ZN => n2332);
   U2388 : OAI22_X1 port map( A1 => n441, A2 => n1864, B1 => n409, B2 => n1865,
                           ZN => n2333);
   U2389 : AOI221_X1 port map( B1 => n1866, B2 => n3964, C1 => n1867, C2 => 
                           n3996, A => n2334, ZN => n2331);
   U2390 : OAI22_X1 port map( A1 => n313, A2 => n1869, B1 => n281, B2 => n1870,
                           ZN => n2334);
   U2391 : AOI221_X1 port map( B1 => n1871, B2 => n177, C1 => n1872, C2 => n49,
                           A => n2335, ZN => n2330);
   U2392 : OAI22_X1 port map( A1 => n113, A2 => n1874, B1 => n241, B2 => n1875,
                           ZN => n2335);
   U2393 : AOI221_X1 port map( B1 => n1876, B2 => n178, C1 => n1877, C2 => n50,
                           A => n2336, ZN => n2329);
   U2394 : OAI22_X1 port map( A1 => n114, A2 => n1879, B1 => n242, B2 => n1880,
                           ZN => n2336);
   U2395 : OAI22_X1 port map( A1 => n2491, A2 => n1828, B1 => n2337, B2 => 
                           n1830, ZN => n2533);
   U2396 : NOR2_X1 port map( A1 => n2338, A2 => n2339, ZN => n2337);
   U2397 : NAND4_X1 port map( A1 => n2340, A2 => n2341, A3 => n2342, A4 => 
                           n2343, ZN => n2339);
   U2398 : AOI221_X1 port map( B1 => n1837, B2 => n3643, C1 => n1838, C2 => 
                           n3675, A => n2344, ZN => n2343);
   U2399 : OAI22_X1 port map( A1 => n1018, A2 => n1840, B1 => n986, B2 => n1841
                           , ZN => n2344);
   U2400 : AOI221_X1 port map( B1 => n1842, B2 => n3707, C1 => n1843, C2 => 
                           n3739, A => n2345, ZN => n2342);
   U2401 : OAI22_X1 port map( A1 => n890, A2 => n1845, B1 => n858, B2 => n1846,
                           ZN => n2345);
   U2402 : AOI221_X1 port map( B1 => n1847, B2 => n3771, C1 => n1848, C2 => 
                           n3803, A => n2346, ZN => n2341);
   U2403 : OAI22_X1 port map( A1 => n698, A2 => n1850, B1 => n666, B2 => n1851,
                           ZN => n2346);
   U2404 : AOI221_X1 port map( B1 => n1852, B2 => n3835, C1 => n1853, C2 => 
                           n3867, A => n2347, ZN => n2340);
   U2405 : OAI22_X1 port map( A1 => n570, A2 => n1855, B1 => n538, B2 => n1856,
                           ZN => n2347);
   U2406 : NAND4_X1 port map( A1 => n2348, A2 => n2349, A3 => n2350, A4 => 
                           n2351, ZN => n2338);
   U2407 : AOI221_X1 port map( B1 => n1861, B2 => n3899, C1 => n1862, C2 => 
                           n3931, A => n2352, ZN => n2351);
   U2408 : OAI22_X1 port map( A1 => n442, A2 => n1864, B1 => n410, B2 => n1865,
                           ZN => n2352);
   U2409 : AOI221_X1 port map( B1 => n1866, B2 => n3963, C1 => n1867, C2 => 
                           n3995, A => n2353, ZN => n2350);
   U2410 : OAI22_X1 port map( A1 => n314, A2 => n1869, B1 => n282, B2 => n1870,
                           ZN => n2353);
   U2411 : AOI221_X1 port map( B1 => n1871, B2 => n179, C1 => n1872, C2 => n51,
                           A => n2354, ZN => n2349);
   U2412 : OAI22_X1 port map( A1 => n115, A2 => n1874, B1 => n243, B2 => n1875,
                           ZN => n2354);
   U2413 : AOI221_X1 port map( B1 => n1876, B2 => n180, C1 => n1877, C2 => n52,
                           A => n2355, ZN => n2348);
   U2414 : OAI22_X1 port map( A1 => n116, A2 => n1879, B1 => n244, B2 => n1880,
                           ZN => n2355);
   U2415 : OAI22_X1 port map( A1 => n2490, A2 => n1828, B1 => n2356, B2 => 
                           n1830, ZN => n2532);
   U2416 : NOR2_X1 port map( A1 => n2357, A2 => n2358, ZN => n2356);
   U2417 : NAND4_X1 port map( A1 => n2359, A2 => n2360, A3 => n2361, A4 => 
                           n2362, ZN => n2358);
   U2418 : AOI221_X1 port map( B1 => n1837, B2 => n3642, C1 => n1838, C2 => 
                           n3674, A => n2363, ZN => n2362);
   U2419 : OAI22_X1 port map( A1 => n1019, A2 => n1840, B1 => n987, B2 => n1841
                           , ZN => n2363);
   U2420 : AOI221_X1 port map( B1 => n1842, B2 => n3706, C1 => n1843, C2 => 
                           n3738, A => n2364, ZN => n2361);
   U2421 : OAI22_X1 port map( A1 => n891, A2 => n1845, B1 => n859, B2 => n1846,
                           ZN => n2364);
   U2422 : AOI221_X1 port map( B1 => n1847, B2 => n3770, C1 => n1848, C2 => 
                           n3802, A => n2365, ZN => n2360);
   U2423 : OAI22_X1 port map( A1 => n699, A2 => n1850, B1 => n667, B2 => n1851,
                           ZN => n2365);
   U2424 : AOI221_X1 port map( B1 => n1852, B2 => n3834, C1 => n1853, C2 => 
                           n3866, A => n2366, ZN => n2359);
   U2425 : OAI22_X1 port map( A1 => n571, A2 => n1855, B1 => n539, B2 => n1856,
                           ZN => n2366);
   U2426 : NAND4_X1 port map( A1 => n2367, A2 => n2368, A3 => n2369, A4 => 
                           n2370, ZN => n2357);
   U2427 : AOI221_X1 port map( B1 => n1861, B2 => n3898, C1 => n1862, C2 => 
                           n3930, A => n2371, ZN => n2370);
   U2428 : OAI22_X1 port map( A1 => n443, A2 => n1864, B1 => n411, B2 => n1865,
                           ZN => n2371);
   U2429 : AOI221_X1 port map( B1 => n1866, B2 => n3962, C1 => n1867, C2 => 
                           n3994, A => n2372, ZN => n2369);
   U2430 : OAI22_X1 port map( A1 => n315, A2 => n1869, B1 => n283, B2 => n1870,
                           ZN => n2372);
   U2431 : AOI221_X1 port map( B1 => n1871, B2 => n181, C1 => n1872, C2 => n53,
                           A => n2373, ZN => n2368);
   U2432 : OAI22_X1 port map( A1 => n117, A2 => n1874, B1 => n245, B2 => n1875,
                           ZN => n2373);
   U2433 : AOI221_X1 port map( B1 => n1876, B2 => n182, C1 => n1877, C2 => n54,
                           A => n2374, ZN => n2367);
   U2434 : OAI22_X1 port map( A1 => n118, A2 => n1879, B1 => n246, B2 => n1880,
                           ZN => n2374);
   U2435 : OAI22_X1 port map( A1 => n2489, A2 => n1828, B1 => n2375, B2 => 
                           n1830, ZN => n2531);
   U2436 : NOR2_X1 port map( A1 => n2376, A2 => n2377, ZN => n2375);
   U2437 : NAND4_X1 port map( A1 => n2378, A2 => n2379, A3 => n2380, A4 => 
                           n2381, ZN => n2377);
   U2438 : AOI221_X1 port map( B1 => n1837, B2 => n3641, C1 => n1838, C2 => 
                           n3673, A => n2382, ZN => n2381);
   U2439 : OAI22_X1 port map( A1 => n1020, A2 => n1840, B1 => n988, B2 => n1841
                           , ZN => n2382);
   U2440 : AOI221_X1 port map( B1 => n1842, B2 => n3705, C1 => n1843, C2 => 
                           n3737, A => n2383, ZN => n2380);
   U2441 : OAI22_X1 port map( A1 => n892, A2 => n1845, B1 => n860, B2 => n1846,
                           ZN => n2383);
   U2442 : AOI221_X1 port map( B1 => n1847, B2 => n3769, C1 => n1848, C2 => 
                           n3801, A => n2384, ZN => n2379);
   U2443 : OAI22_X1 port map( A1 => n700, A2 => n1850, B1 => n668, B2 => n1851,
                           ZN => n2384);
   U2444 : AOI221_X1 port map( B1 => n1852, B2 => n3833, C1 => n1853, C2 => 
                           n3865, A => n2385, ZN => n2378);
   U2445 : OAI22_X1 port map( A1 => n572, A2 => n1855, B1 => n540, B2 => n1856,
                           ZN => n2385);
   U2446 : NAND4_X1 port map( A1 => n2386, A2 => n2387, A3 => n2388, A4 => 
                           n2389, ZN => n2376);
   U2447 : AOI221_X1 port map( B1 => n1861, B2 => n3897, C1 => n1862, C2 => 
                           n3929, A => n2390, ZN => n2389);
   U2448 : OAI22_X1 port map( A1 => n444, A2 => n1864, B1 => n412, B2 => n1865,
                           ZN => n2390);
   U2449 : AOI221_X1 port map( B1 => n1866, B2 => n3961, C1 => n1867, C2 => 
                           n3993, A => n2391, ZN => n2388);
   U2450 : OAI22_X1 port map( A1 => n316, A2 => n1869, B1 => n284, B2 => n1870,
                           ZN => n2391);
   U2451 : AOI221_X1 port map( B1 => n1871, B2 => n183, C1 => n1872, C2 => n55,
                           A => n2392, ZN => n2387);
   U2452 : OAI22_X1 port map( A1 => n119, A2 => n1874, B1 => n247, B2 => n1875,
                           ZN => n2392);
   U2453 : AOI221_X1 port map( B1 => n1876, B2 => n184, C1 => n1877, C2 => n56,
                           A => n2393, ZN => n2386);
   U2454 : OAI22_X1 port map( A1 => n120, A2 => n1879, B1 => n248, B2 => n1880,
                           ZN => n2393);
   U2455 : OAI22_X1 port map( A1 => n2488, A2 => n1828, B1 => n2394, B2 => 
                           n1830, ZN => n2530);
   U2456 : NOR2_X1 port map( A1 => n2395, A2 => n2396, ZN => n2394);
   U2457 : NAND4_X1 port map( A1 => n2397, A2 => n2398, A3 => n2399, A4 => 
                           n2400, ZN => n2396);
   U2458 : AOI221_X1 port map( B1 => n1837, B2 => n3640, C1 => n1838, C2 => 
                           n3672, A => n2401, ZN => n2400);
   U2459 : OAI22_X1 port map( A1 => n1021, A2 => n1840, B1 => n989, B2 => n1841
                           , ZN => n2401);
   U2460 : AOI221_X1 port map( B1 => n1842, B2 => n3704, C1 => n1843, C2 => 
                           n3736, A => n2402, ZN => n2399);
   U2461 : OAI22_X1 port map( A1 => n893, A2 => n1845, B1 => n861, B2 => n1846,
                           ZN => n2402);
   U2462 : AOI221_X1 port map( B1 => n1847, B2 => n3768, C1 => n1848, C2 => 
                           n3800, A => n2403, ZN => n2398);
   U2463 : OAI22_X1 port map( A1 => n701, A2 => n1850, B1 => n669, B2 => n1851,
                           ZN => n2403);
   U2464 : AOI221_X1 port map( B1 => n1852, B2 => n3832, C1 => n1853, C2 => 
                           n3864, A => n2404, ZN => n2397);
   U2465 : OAI22_X1 port map( A1 => n573, A2 => n1855, B1 => n541, B2 => n1856,
                           ZN => n2404);
   U2466 : NAND4_X1 port map( A1 => n2405, A2 => n2406, A3 => n2407, A4 => 
                           n2408, ZN => n2395);
   U2467 : AOI221_X1 port map( B1 => n1861, B2 => n3896, C1 => n1862, C2 => 
                           n3928, A => n2409, ZN => n2408);
   U2468 : OAI22_X1 port map( A1 => n445, A2 => n1864, B1 => n413, B2 => n1865,
                           ZN => n2409);
   U2469 : AOI221_X1 port map( B1 => n1866, B2 => n3960, C1 => n1867, C2 => 
                           n3992, A => n2410, ZN => n2407);
   U2470 : OAI22_X1 port map( A1 => n317, A2 => n1869, B1 => n285, B2 => n1870,
                           ZN => n2410);
   U2471 : AOI221_X1 port map( B1 => n1871, B2 => n185, C1 => n1872, C2 => n57,
                           A => n2411, ZN => n2406);
   U2472 : OAI22_X1 port map( A1 => n121, A2 => n1874, B1 => n249, B2 => n1875,
                           ZN => n2411);
   U2473 : AOI221_X1 port map( B1 => n1876, B2 => n186, C1 => n1877, C2 => n58,
                           A => n2412, ZN => n2405);
   U2474 : OAI22_X1 port map( A1 => n122, A2 => n1879, B1 => n250, B2 => n1880,
                           ZN => n2412);
   U2475 : OAI22_X1 port map( A1 => n2487, A2 => n1828, B1 => n2413, B2 => 
                           n1830, ZN => n2529);
   U2476 : NOR2_X1 port map( A1 => n2414, A2 => n2415, ZN => n2413);
   U2477 : NAND4_X1 port map( A1 => n2416, A2 => n2417, A3 => n2418, A4 => 
                           n2419, ZN => n2415);
   U2478 : AOI221_X1 port map( B1 => n1837, B2 => n3639, C1 => n1838, C2 => 
                           n3671, A => n2420, ZN => n2419);
   U2479 : OAI22_X1 port map( A1 => n1022, A2 => n1840, B1 => n990, B2 => n1841
                           , ZN => n2420);
   U2480 : AOI221_X1 port map( B1 => n1842, B2 => n3703, C1 => n1843, C2 => 
                           n3735, A => n2421, ZN => n2418);
   U2481 : OAI22_X1 port map( A1 => n894, A2 => n1845, B1 => n862, B2 => n1846,
                           ZN => n2421);
   U2482 : AOI221_X1 port map( B1 => n1847, B2 => n3767, C1 => n1848, C2 => 
                           n3799, A => n2422, ZN => n2417);
   U2483 : OAI22_X1 port map( A1 => n702, A2 => n1850, B1 => n670, B2 => n1851,
                           ZN => n2422);
   U2484 : AOI221_X1 port map( B1 => n1852, B2 => n3831, C1 => n1853, C2 => 
                           n3863, A => n2423, ZN => n2416);
   U2485 : OAI22_X1 port map( A1 => n574, A2 => n1855, B1 => n542, B2 => n1856,
                           ZN => n2423);
   U2486 : NAND4_X1 port map( A1 => n2424, A2 => n2425, A3 => n2426, A4 => 
                           n2427, ZN => n2414);
   U2487 : AOI221_X1 port map( B1 => n1861, B2 => n3895, C1 => n1862, C2 => 
                           n3927, A => n2428, ZN => n2427);
   U2488 : OAI22_X1 port map( A1 => n446, A2 => n1864, B1 => n414, B2 => n1865,
                           ZN => n2428);
   U2489 : AOI221_X1 port map( B1 => n1866, B2 => n3959, C1 => n1867, C2 => 
                           n3991, A => n2429, ZN => n2426);
   U2490 : OAI22_X1 port map( A1 => n318, A2 => n1869, B1 => n286, B2 => n1870,
                           ZN => n2429);
   U2491 : AOI221_X1 port map( B1 => n1871, B2 => n187, C1 => n1872, C2 => n59,
                           A => n2430, ZN => n2425);
   U2492 : OAI22_X1 port map( A1 => n123, A2 => n1874, B1 => n251, B2 => n1875,
                           ZN => n2430);
   U2493 : AOI221_X1 port map( B1 => n1876, B2 => n188, C1 => n1877, C2 => n60,
                           A => n2431, ZN => n2424);
   U2494 : OAI22_X1 port map( A1 => n124, A2 => n1879, B1 => n252, B2 => n1880,
                           ZN => n2431);
   U2495 : OAI22_X1 port map( A1 => n2486, A2 => n1828, B1 => n2432, B2 => 
                           n1830, ZN => n2528);
   U2496 : NOR2_X1 port map( A1 => n2433, A2 => n2434, ZN => n2432);
   U2497 : NAND4_X1 port map( A1 => n2435, A2 => n2436, A3 => n2437, A4 => 
                           n2438, ZN => n2434);
   U2498 : AOI221_X1 port map( B1 => n1837, B2 => n3638, C1 => n1838, C2 => 
                           n3670, A => n2439, ZN => n2438);
   U2499 : OAI22_X1 port map( A1 => n1023, A2 => n1840, B1 => n991, B2 => n1841
                           , ZN => n2439);
   U2500 : AOI221_X1 port map( B1 => n1842, B2 => n3702, C1 => n1843, C2 => 
                           n3734, A => n2440, ZN => n2437);
   U2501 : OAI22_X1 port map( A1 => n895, A2 => n1845, B1 => n863, B2 => n1846,
                           ZN => n2440);
   U2502 : AOI221_X1 port map( B1 => n1847, B2 => n3766, C1 => n1848, C2 => 
                           n3798, A => n2441, ZN => n2436);
   U2503 : OAI22_X1 port map( A1 => n703, A2 => n1850, B1 => n671, B2 => n1851,
                           ZN => n2441);
   U2504 : AOI221_X1 port map( B1 => n1852, B2 => n3830, C1 => n1853, C2 => 
                           n3862, A => n2442, ZN => n2435);
   U2505 : OAI22_X1 port map( A1 => n575, A2 => n1855, B1 => n543, B2 => n1856,
                           ZN => n2442);
   U2506 : NAND4_X1 port map( A1 => n2443, A2 => n2444, A3 => n2445, A4 => 
                           n2446, ZN => n2433);
   U2507 : AOI221_X1 port map( B1 => n1861, B2 => n3894, C1 => n1862, C2 => 
                           n3926, A => n2447, ZN => n2446);
   U2508 : OAI22_X1 port map( A1 => n447, A2 => n1864, B1 => n415, B2 => n1865,
                           ZN => n2447);
   U2509 : AOI221_X1 port map( B1 => n1866, B2 => n3958, C1 => n1867, C2 => 
                           n3990, A => n2448, ZN => n2445);
   U2510 : OAI22_X1 port map( A1 => n319, A2 => n1869, B1 => n287, B2 => n1870,
                           ZN => n2448);
   U2511 : AOI221_X1 port map( B1 => n1871, B2 => n189, C1 => n1872, C2 => n61,
                           A => n2449, ZN => n2444);
   U2512 : OAI22_X1 port map( A1 => n125, A2 => n1874, B1 => n253, B2 => n1875,
                           ZN => n2449);
   U2513 : AOI221_X1 port map( B1 => n1876, B2 => n190, C1 => n1877, C2 => n62,
                           A => n2450, ZN => n2443);
   U2514 : OAI22_X1 port map( A1 => n126, A2 => n1879, B1 => n254, B2 => n1880,
                           ZN => n2450);
   U2515 : OAI22_X1 port map( A1 => n2485, A2 => n1828, B1 => n2451, B2 => 
                           n1830, ZN => n2527);
   U2516 : NOR2_X1 port map( A1 => n2452, A2 => n2453, ZN => n2451);
   U2517 : NAND4_X1 port map( A1 => n2454, A2 => n2455, A3 => n2456, A4 => 
                           n2457, ZN => n2453);
   U2518 : AOI221_X1 port map( B1 => n1837, B2 => n3637, C1 => n1838, C2 => 
                           n3669, A => n2458, ZN => n2457);
   U2519 : OAI22_X1 port map( A1 => n1024, A2 => n1840, B1 => n992, B2 => n1841
                           , ZN => n2458);
   U2520 : AOI221_X1 port map( B1 => n1842, B2 => n3701, C1 => n1843, C2 => 
                           n3733, A => n2463, ZN => n2456);
   U2521 : OAI22_X1 port map( A1 => n896, A2 => n1845, B1 => n864, B2 => n1846,
                           ZN => n2463);
   U2522 : AND3_X1 port map( A1 => ADD_RD2(3), A2 => n2466, A3 => ADD_RD2(4), 
                           ZN => n2459);
   U2523 : AND3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(0), A3 => 
                           ADD_RD2(4), ZN => n2461);
   U2524 : AOI221_X1 port map( B1 => n1847, B2 => n3765, C1 => n1848, C2 => 
                           n3797, A => n2467, ZN => n2455);
   U2525 : OAI22_X1 port map( A1 => n704, A2 => n1850, B1 => n672, B2 => n1851,
                           ZN => n2467);
   U2526 : AOI221_X1 port map( B1 => n1852, B2 => n3829, C1 => n1853, C2 => 
                           n3861, A => n2470, ZN => n2454);
   U2527 : OAI22_X1 port map( A1 => n576, A2 => n1855, B1 => n544, B2 => n1856,
                           ZN => n2470);
   U2528 : AND3_X1 port map( A1 => n2466, A2 => n2471, A3 => ADD_RD2(4), ZN => 
                           n2468);
   U2529 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => n2471, A3 => ADD_RD2(4), 
                           ZN => n2469);
   U2530 : NAND4_X1 port map( A1 => n2472, A2 => n2473, A3 => n2474, A4 => 
                           n2475, ZN => n2452);
   U2531 : AOI221_X1 port map( B1 => n1861, B2 => n3893, C1 => n1862, C2 => 
                           n3925, A => n2476, ZN => n2475);
   U2532 : OAI22_X1 port map( A1 => n448, A2 => n1864, B1 => n416, B2 => n1865,
                           ZN => n2476);
   U2533 : AOI221_X1 port map( B1 => n1866, B2 => n3957, C1 => n1867, C2 => 
                           n3989, A => n2479, ZN => n2474);
   U2534 : OAI22_X1 port map( A1 => n320, A2 => n1869, B1 => n288, B2 => n1870,
                           ZN => n2479);
   U2535 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n2471, 
                           ZN => n2477);
   U2536 : NOR3_X1 port map( A1 => n2466, A2 => ADD_RD2(4), A3 => n2471, ZN => 
                           n2478);
   U2537 : INV_X1 port map( A => ADD_RD2(3), ZN => n2471);
   U2538 : AOI221_X1 port map( B1 => n1871, B2 => n191, C1 => n1872, C2 => n63,
                           A => n2480, ZN => n2473);
   U2539 : OAI22_X1 port map( A1 => n127, A2 => n1874, B1 => n255, B2 => n1875,
                           ZN => n2480);
   U2540 : AND2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), ZN => n2460);
   U2541 : AND2_X1 port map( A1 => ADD_RD2(2), A2 => n2483, ZN => n2462);
   U2542 : AOI221_X1 port map( B1 => n1876, B2 => n192, C1 => n1877, C2 => n64,
                           A => n2484, ZN => n2472);
   U2543 : OAI22_X1 port map( A1 => n128, A2 => n1879, B1 => n256, B2 => n1880,
                           ZN => n2484);
   U2544 : NOR2_X1 port map( A1 => n2483, A2 => ADD_RD2(2), ZN => n2464);
   U2545 : INV_X1 port map( A => ADD_RD2(1), ZN => n2483);
   U2546 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n2466, 
                           ZN => n2481);
   U2547 : INV_X1 port map( A => ADD_RD2(0), ZN => n2466);
   U2548 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n2465);
   U2549 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n2482);
   U2550 : INV_X1 port map( A => RST, ZN => n1827);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ADDER_N32 is

   port( CURR_ADDR : in std_logic_vector (31 downto 0);  NEXT_ADDR : out 
         std_logic_vector (31 downto 0));

end ADDER_N32;

architecture SYN_BEHAVIOR of ADDER_N32 is

   component ADDER_N32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n3, n_1556 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '1';
   n3 <= '0';
   add_26 : ADDER_N32_DW01_add_0 port map( A(31) => CURR_ADDR(31), A(30) => 
                           CURR_ADDR(30), A(29) => CURR_ADDR(29), A(28) => 
                           CURR_ADDR(28), A(27) => CURR_ADDR(27), A(26) => 
                           CURR_ADDR(26), A(25) => CURR_ADDR(25), A(24) => 
                           CURR_ADDR(24), A(23) => CURR_ADDR(23), A(22) => 
                           CURR_ADDR(22), A(21) => CURR_ADDR(21), A(20) => 
                           CURR_ADDR(20), A(19) => CURR_ADDR(19), A(18) => 
                           CURR_ADDR(18), A(17) => CURR_ADDR(17), A(16) => 
                           CURR_ADDR(16), A(15) => CURR_ADDR(15), A(14) => 
                           CURR_ADDR(14), A(13) => CURR_ADDR(13), A(12) => 
                           CURR_ADDR(12), A(11) => CURR_ADDR(11), A(10) => 
                           CURR_ADDR(10), A(9) => CURR_ADDR(9), A(8) => 
                           CURR_ADDR(8), A(7) => CURR_ADDR(7), A(6) => 
                           CURR_ADDR(6), A(5) => CURR_ADDR(5), A(4) => 
                           CURR_ADDR(4), A(3) => CURR_ADDR(3), A(2) => 
                           CURR_ADDR(2), A(1) => CURR_ADDR(1), A(0) => 
                           CURR_ADDR(0), B(31) => n1, B(30) => n1, B(29) => n1,
                           B(28) => n1, B(27) => n1, B(26) => n1, B(25) => n1, 
                           B(24) => n1, B(23) => n1, B(22) => n1, B(21) => n1, 
                           B(20) => n1, B(19) => n1, B(18) => n1, B(17) => n1, 
                           B(16) => n1, B(15) => n1, B(14) => n1, B(13) => n1, 
                           B(12) => n1, B(11) => n1, B(10) => n1, B(9) => n1, 
                           B(8) => n1, B(7) => n1, B(6) => n1, B(5) => n1, B(4)
                           => n1, B(3) => n1, B(2) => n2, B(1) => n1, B(0) => 
                           n1, CI => n3, SUM(31) => NEXT_ADDR(31), SUM(30) => 
                           NEXT_ADDR(30), SUM(29) => NEXT_ADDR(29), SUM(28) => 
                           NEXT_ADDR(28), SUM(27) => NEXT_ADDR(27), SUM(26) => 
                           NEXT_ADDR(26), SUM(25) => NEXT_ADDR(25), SUM(24) => 
                           NEXT_ADDR(24), SUM(23) => NEXT_ADDR(23), SUM(22) => 
                           NEXT_ADDR(22), SUM(21) => NEXT_ADDR(21), SUM(20) => 
                           NEXT_ADDR(20), SUM(19) => NEXT_ADDR(19), SUM(18) => 
                           NEXT_ADDR(18), SUM(17) => NEXT_ADDR(17), SUM(16) => 
                           NEXT_ADDR(16), SUM(15) => NEXT_ADDR(15), SUM(14) => 
                           NEXT_ADDR(14), SUM(13) => NEXT_ADDR(13), SUM(12) => 
                           NEXT_ADDR(12), SUM(11) => NEXT_ADDR(11), SUM(10) => 
                           NEXT_ADDR(10), SUM(9) => NEXT_ADDR(9), SUM(8) => 
                           NEXT_ADDR(8), SUM(7) => NEXT_ADDR(7), SUM(6) => 
                           NEXT_ADDR(6), SUM(5) => NEXT_ADDR(5), SUM(4) => 
                           NEXT_ADDR(4), SUM(3) => NEXT_ADDR(3), SUM(2) => 
                           NEXT_ADDR(2), SUM(1) => NEXT_ADDR(1), SUM(0) => 
                           NEXT_ADDR(0), CO => n_1556);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT5_0 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_GENERIC_NBIT5_0;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT5_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U5 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21 is

   port( A, B, SEL : in std_logic;  Y : out std_logic);

end MUX21;

architecture SYN_BEHAVIOR of MUX21 is

   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X2 port map( A => A, B => B, S => SEL, Z => Y);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_GENERIC_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_0;

architecture SYN_BEHAVIOR of MUX21_GENERIC_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BRANCHING_UNIT_N32 is

   port( CLK, RST : in std_logic;  Reg_A : in std_logic_vector (31 downto 0);  
         EQ_cond, IS_JUMP : in std_logic;  branch_taken : out std_logic);

end BRANCHING_UNIT_N32;

architecture SYN_BEHAVIOR of BRANCHING_UNIT_N32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n_1557 :
      std_logic;

begin
   
   branch_taken_reg : DFF_X1 port map( D => n14, CK => CLK, Q => branch_taken, 
                           QN => n_1557);
   U3 : INV_X1 port map( A => n1, ZN => n14);
   U4 : OAI21_X1 port map( B1 => IS_JUMP, B2 => n2, A => RST, ZN => n1);
   U5 : XNOR2_X1 port map( A => EQ_cond, B => n3, ZN => n2);
   U6 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n3);
   U7 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n5);
   U8 : NOR4_X1 port map( A1 => Reg_A(23), A2 => Reg_A(22), A3 => Reg_A(21), A4
                           => Reg_A(20), ZN => n9);
   U9 : NOR4_X1 port map( A1 => Reg_A(1), A2 => Reg_A(19), A3 => Reg_A(18), A4 
                           => Reg_A(17), ZN => n8);
   U10 : NOR4_X1 port map( A1 => Reg_A(16), A2 => Reg_A(15), A3 => Reg_A(14), 
                           A4 => Reg_A(13), ZN => n7);
   U11 : NOR4_X1 port map( A1 => Reg_A(12), A2 => Reg_A(11), A3 => Reg_A(10), 
                           A4 => Reg_A(0), ZN => n6);
   U12 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12, A4 => n13, ZN => 
                           n4);
   U13 : NOR4_X1 port map( A1 => Reg_A(9), A2 => Reg_A(8), A3 => Reg_A(7), A4 
                           => Reg_A(6), ZN => n13);
   U14 : NOR4_X1 port map( A1 => Reg_A(5), A2 => Reg_A(4), A3 => Reg_A(3), A4 
                           => Reg_A(31), ZN => n12);
   U15 : NOR4_X1 port map( A1 => Reg_A(30), A2 => Reg_A(2), A3 => Reg_A(29), A4
                           => Reg_A(28), ZN => n11);
   U16 : NOR4_X1 port map( A1 => Reg_A(27), A2 => Reg_A(26), A3 => Reg_A(25), 
                           A4 => Reg_A(24), ZN => n10);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT5_0 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 downto 
         0);  DATA_OUT : out std_logic_vector (4 downto 0));

end REG_GENERIC_NBIT5_0;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n14, CK => CLK, Q => DATA_OUT(4)
                           , QN => n13);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n15, CK => CLK, Q => DATA_OUT(3)
                           , QN => n12);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n16, CK => CLK, Q => DATA_OUT(2)
                           , QN => n11);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n17, CK => CLK, Q => DATA_OUT(1)
                           , QN => n10);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n18, CK => CLK, Q => DATA_OUT(0)
                           , QN => n9);
   U3 : OAI21_X1 port map( B1 => n13, B2 => n1, A => n2, ZN => n14);
   U4 : NAND2_X1 port map( A1 => DATA_IN(4), A2 => n3, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n12, B2 => n1, A => n4, ZN => n15);
   U6 : NAND2_X1 port map( A1 => DATA_IN(3), A2 => n3, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n11, B2 => n1, A => n5, ZN => n16);
   U8 : NAND2_X1 port map( A1 => DATA_IN(2), A2 => n3, ZN => n5);
   U9 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n6, ZN => n17);
   U10 : NAND2_X1 port map( A1 => DATA_IN(1), A2 => n3, ZN => n6);
   U11 : OAI21_X1 port map( B1 => n9, B2 => n1, A => n7, ZN => n18);
   U12 : NAND2_X1 port map( A1 => DATA_IN(0), A2 => n3, ZN => n7);
   U13 : AND2_X1 port map( A1 => RST, A2 => n1, ZN => n3);
   U14 : NAND2_X1 port map( A1 => n8, A2 => RST, ZN => n1);
   U15 : INV_X1 port map( A => EN, ZN => n8);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT26 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (25 downto
         0);  DATA_OUT : out std_logic_vector (25 downto 0));

end REG_GENERIC_NBIT26;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81 : std_logic;

begin
   
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n56, CK => CLK, Q => 
                           DATA_OUT(25), QN => n55);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n57, CK => CLK, Q => 
                           DATA_OUT(24), QN => n54);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n58, CK => CLK, Q => 
                           DATA_OUT(23), QN => n53);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n59, CK => CLK, Q => 
                           DATA_OUT(22), QN => n52);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n60, CK => CLK, Q => 
                           DATA_OUT(21), QN => n51);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n61, CK => CLK, Q => 
                           DATA_OUT(20), QN => n50);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n62, CK => CLK, Q => 
                           DATA_OUT(19), QN => n49);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n63, CK => CLK, Q => 
                           DATA_OUT(18), QN => n48);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n64, CK => CLK, Q => 
                           DATA_OUT(17), QN => n47);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n65, CK => CLK, Q => 
                           DATA_OUT(16), QN => n46);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n66, CK => CLK, Q => 
                           DATA_OUT(15), QN => n45);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n67, CK => CLK, Q => 
                           DATA_OUT(14), QN => n44);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(13), QN => n43);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(12), QN => n42);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(11), QN => n41);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(10), QN => n40);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n72, CK => CLK, Q => DATA_OUT(9)
                           , QN => n39);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n73, CK => CLK, Q => DATA_OUT(8)
                           , QN => n38);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n74, CK => CLK, Q => DATA_OUT(7)
                           , QN => n37);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n75, CK => CLK, Q => DATA_OUT(6)
                           , QN => n36);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n76, CK => CLK, Q => DATA_OUT(5)
                           , QN => n35);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n77, CK => CLK, Q => DATA_OUT(4)
                           , QN => n34);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n78, CK => CLK, Q => DATA_OUT(3)
                           , QN => n33);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n79, CK => CLK, Q => DATA_OUT(2)
                           , QN => n32);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n80, CK => CLK, Q => DATA_OUT(1)
                           , QN => n31);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n81, CK => CLK, Q => DATA_OUT(0)
                           , QN => n30);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n29, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n3, ZN => n56);
   U6 : INV_X1 port map( A => DATA_IN(25), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n4, ZN => n57);
   U8 : INV_X1 port map( A => DATA_IN(24), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n5, ZN => n58);
   U10 : INV_X1 port map( A => DATA_IN(23), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n6, ZN => n59)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(22), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n7, ZN => n60)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(21), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n8, ZN => n61)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(20), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n9, ZN => n62)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(19), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n10, ZN => n63
                           );
   U20 : INV_X1 port map( A => DATA_IN(18), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n11, ZN => n64
                           );
   U22 : INV_X1 port map( A => DATA_IN(17), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n12, ZN => n65
                           );
   U24 : INV_X1 port map( A => DATA_IN(16), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n13, ZN => n66
                           );
   U26 : INV_X1 port map( A => DATA_IN(15), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n14, ZN => n67
                           );
   U28 : INV_X1 port map( A => DATA_IN(14), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n15, ZN => n68
                           );
   U30 : INV_X1 port map( A => DATA_IN(13), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n16, ZN => n69
                           );
   U32 : INV_X1 port map( A => DATA_IN(12), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n17, ZN => n70
                           );
   U34 : INV_X1 port map( A => DATA_IN(11), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n18, ZN => n71
                           );
   U36 : INV_X1 port map( A => DATA_IN(10), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n19, ZN => n72
                           );
   U38 : INV_X1 port map( A => DATA_IN(9), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n20, ZN => n73
                           );
   U40 : INV_X1 port map( A => DATA_IN(8), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n21, ZN => n74
                           );
   U42 : INV_X1 port map( A => DATA_IN(7), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n22, ZN => n75
                           );
   U44 : INV_X1 port map( A => DATA_IN(6), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n35, A2 => n1, B1 => n2, B2 => n23, ZN => n76
                           );
   U46 : INV_X1 port map( A => DATA_IN(5), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n34, A2 => n1, B1 => n2, B2 => n24, ZN => n77
                           );
   U48 : INV_X1 port map( A => DATA_IN(4), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n33, A2 => n1, B1 => n2, B2 => n25, ZN => n78
                           );
   U50 : INV_X1 port map( A => DATA_IN(3), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n32, A2 => n1, B1 => n2, B2 => n26, ZN => n79
                           );
   U52 : INV_X1 port map( A => DATA_IN(2), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n31, A2 => n1, B1 => n2, B2 => n27, ZN => n80
                           );
   U54 : INV_X1 port map( A => DATA_IN(1), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n30, A2 => n1, B1 => n2, B2 => n28, ZN => n81
                           );
   U56 : INV_X1 port map( A => DATA_IN(0), ZN => n28);
   U57 : INV_X1 port map( A => EN, ZN => n29);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity dlx_cu is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
         EQ_COND, IS_JUMP : out std_logic;  ALU_OPCODE : out std_logic_vector 
         (0 to 3);  DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, IS_JAL, 
         WB_MUX_SEL, RF_WE : out std_logic);

end dlx_cu;

architecture SYN_dlx_cu_hw of dlx_cu is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal cw_17_port, cw_14_port, cw_13_port, cw_12_port, cw_9_port, cw_8_port,
      cw_6_port, cw_5_port, cw_4_port, cw_3_port, cw_1_port, cw2_12_port, 
      cw2_11_port, cw2_10_port, cw2_9_port, cw2_8_port, cw2_7_port, cw2_6_port,
      cw2_5_port, cw2_4_port, cw2_3_port, cw2_2_port, cw2_1_port, cw2_0_port, 
      cw3_6_port, cw3_5_port, cw3_4_port, cw3_3_port, cw3_2_port, cw3_1_port, 
      cw3_0_port, cw4_2_port, cw4_1_port, cw4_0_port, aluOpcode1_3_port, 
      aluOpcode1_2_port, aluOpcode1_1_port, aluOpcode1_0_port, 
      aluOpcode_i_3_port, aluOpcode_i_2_port, aluOpcode_i_1_port, 
      aluOpcode_i_0_port, n1, n2, n34, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606 : std_logic;

begin
   
   cw2_reg_15_inst : DFFR_X1 port map( D => cw_9_port, CK => Clk, RN => Rst, Q 
                           => RegA_LATCH_EN, QN => n_1558);
   cw2_reg_14_inst : DFFR_X1 port map( D => cw_14_port, CK => Clk, RN => Rst, Q
                           => RegB_LATCH_EN, QN => n_1559);
   cw2_reg_13_inst : DFFR_X1 port map( D => cw_13_port, CK => Clk, RN => Rst, Q
                           => RegIMM_LATCH_EN, QN => n_1560);
   cw2_reg_12_inst : DFFR_X1 port map( D => cw_12_port, CK => Clk, RN => Rst, Q
                           => cw2_12_port, QN => n_1561);
   cw2_reg_11_inst : DFFR_X1 port map( D => cw_4_port, CK => Clk, RN => Rst, Q 
                           => cw2_11_port, QN => n_1562);
   cw2_reg_10_inst : DFFR_X1 port map( D => cw_13_port, CK => Clk, RN => Rst, Q
                           => cw2_10_port, QN => n_1563);
   cw2_reg_9_inst : DFFR_X1 port map( D => cw_9_port, CK => Clk, RN => Rst, Q 
                           => cw2_9_port, QN => n_1564);
   cw2_reg_8_inst : DFFR_X1 port map( D => cw_8_port, CK => Clk, RN => Rst, Q 
                           => cw2_8_port, QN => n_1565);
   cw2_reg_7_inst : DFFR_X1 port map( D => n66, CK => Clk, RN => Rst, Q => 
                           cw2_7_port, QN => n_1566);
   cw2_reg_6_inst : DFFR_X1 port map( D => cw_6_port, CK => Clk, RN => Rst, Q 
                           => cw2_6_port, QN => n_1567);
   cw2_reg_5_inst : DFFR_X1 port map( D => cw_5_port, CK => Clk, RN => Rst, Q 
                           => cw2_5_port, QN => n_1568);
   cw2_reg_4_inst : DFFR_X1 port map( D => cw_4_port, CK => Clk, RN => Rst, Q 
                           => cw2_4_port, QN => n_1569);
   cw2_reg_3_inst : DFFR_X1 port map( D => cw_3_port, CK => Clk, RN => Rst, Q 
                           => cw2_3_port, QN => n_1570);
   cw2_reg_2_inst : SDFFR_X1 port map( D => n2, SI => n66, SE => IR_IN(26), CK 
                           => Clk, RN => Rst, Q => cw2_2_port, QN => n_1571);
   cw2_reg_1_inst : DFFR_X1 port map( D => cw_1_port, CK => Clk, RN => Rst, Q 
                           => cw2_1_port, QN => n_1572);
   cw2_reg_0_inst : SDFFR_X1 port map( D => n1, SI => cw_1_port, SE => n34, CK 
                           => Clk, RN => Rst, Q => cw2_0_port, QN => n_1573);
   cw1_reg_17_inst : DFFR_X1 port map( D => cw_17_port, CK => Clk, RN => Rst, Q
                           => IR_LATCH_EN, QN => n_1574);
   cw1_reg_16_inst : DFFR_X1 port map( D => cw_17_port, CK => Clk, RN => Rst, Q
                           => NPC_LATCH_EN, QN => n_1575);
   cw3_reg_12_inst : DFFR_X1 port map( D => cw2_12_port, CK => Clk, RN => Rst, 
                           Q => SIGNED_IMM, QN => n_1576);
   cw3_reg_9_inst : DFFR_X1 port map( D => cw2_9_port, CK => Clk, RN => Rst, Q 
                           => ALU_OUTREG_EN, QN => n_1577);
   cw3_reg_8_inst : DFFR_X1 port map( D => cw2_8_port, CK => Clk, RN => Rst, Q 
                           => EQ_COND, QN => n_1578);
   cw3_reg_7_inst : DFFR_X1 port map( D => cw2_7_port, CK => Clk, RN => Rst, Q 
                           => IS_JUMP, QN => n_1579);
   cw3_reg_6_inst : DFFR_X1 port map( D => cw2_6_port, CK => Clk, RN => Rst, Q 
                           => cw3_6_port, QN => n_1580);
   cw3_reg_5_inst : DFFR_X1 port map( D => cw2_5_port, CK => Clk, RN => Rst, Q 
                           => cw3_5_port, QN => n_1581);
   cw3_reg_4_inst : DFFR_X1 port map( D => cw2_4_port, CK => Clk, RN => Rst, Q 
                           => cw3_4_port, QN => n_1582);
   cw3_reg_3_inst : DFFR_X1 port map( D => cw2_3_port, CK => Clk, RN => Rst, Q 
                           => cw3_3_port, QN => n_1583);
   cw3_reg_2_inst : DFFR_X1 port map( D => cw2_2_port, CK => Clk, RN => Rst, Q 
                           => cw3_2_port, QN => n_1584);
   cw3_reg_1_inst : DFFR_X1 port map( D => cw2_1_port, CK => Clk, RN => Rst, Q 
                           => cw3_1_port, QN => n_1585);
   cw3_reg_0_inst : DFFR_X1 port map( D => cw2_0_port, CK => Clk, RN => Rst, Q 
                           => cw3_0_port, QN => n_1586);
   cw4_reg_6_inst : DFFR_X1 port map( D => cw3_6_port, CK => Clk, RN => Rst, Q 
                           => DRAM_WE, QN => n_1587);
   cw4_reg_5_inst : DFFR_X1 port map( D => cw3_5_port, CK => Clk, RN => Rst, Q 
                           => LMD_LATCH_EN, QN => n_1588);
   cw4_reg_4_inst : DFFR_X1 port map( D => cw3_4_port, CK => Clk, RN => Rst, Q 
                           => JUMP_EN, QN => n_1589);
   cw4_reg_2_inst : DFFR_X1 port map( D => cw3_2_port, CK => Clk, RN => Rst, Q 
                           => cw4_2_port, QN => n_1590);
   cw4_reg_1_inst : DFFR_X1 port map( D => cw3_1_port, CK => Clk, RN => Rst, Q 
                           => cw4_1_port, QN => n_1591);
   cw4_reg_0_inst : DFFR_X1 port map( D => cw3_0_port, CK => Clk, RN => Rst, Q 
                           => cw4_0_port, QN => n_1592);
   cw5_reg_0_inst : DFFR_X1 port map( D => cw4_0_port, CK => Clk, RN => Rst, Q 
                           => RF_WE, QN => n_1593);
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_3_port, QN => n_1594);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_2_port, QN => n_1595);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_1_port, QN => n_1596);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_0_port, QN => n_1597);
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => aluOpcode1_3_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(0), QN => n_1598);
   aluOpcode2_reg_2_inst : DFFR_X1 port map( D => aluOpcode1_2_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(1), QN => n_1599);
   aluOpcode2_reg_1_inst : DFFR_X1 port map( D => aluOpcode1_1_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(2), QN => n_1600);
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => aluOpcode1_0_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(3), QN => n_1601);
   n1 <= '1';
   n2 <= '0';
   cw5_reg_2_inst : DFFR_X2 port map( D => cw4_2_port, CK => Clk, RN => Rst, Q 
                           => IS_JAL, QN => n_1602);
   cw3_reg_11_inst : DFFR_X2 port map( D => cw2_11_port, CK => Clk, RN => Rst, 
                           Q => MUXA_SEL, QN => n_1603);
   cw3_reg_10_inst : DFFR_X2 port map( D => cw2_10_port, CK => Clk, RN => Rst, 
                           Q => MUXB_SEL, QN => n_1604);
   cw5_reg_1_inst : DFFR_X2 port map( D => cw4_1_port, CK => Clk, RN => Rst, Q 
                           => WB_MUX_SEL, QN => n_1605);
   cw4_reg_3_inst : DFFR_X2 port map( D => cw3_3_port, CK => Clk, RN => Rst, Q 
                           => PC_LATCH_EN, QN => n_1606);
   U5 : OAI21_X1 port map( B1 => n3, B2 => n4, A => n5, ZN => cw_9_port);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n6, A => n7, ZN => cw_8_port);
   U7 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => n6);
   U8 : NOR2_X1 port map( A1 => IR_IN(29), A2 => n10, ZN => cw_5_port);
   U9 : INV_X1 port map( A => n11, ZN => cw_4_port);
   U10 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => cw_3_port);
   U11 : AND4_X1 port map( A1 => n12, A2 => n13, A3 => n10, A4 => n34, ZN => n5
                           );
   U12 : NAND3_X1 port map( A1 => n14, A2 => n8, A3 => IR_IN(26), ZN => n34);
   U13 : OAI211_X1 port map( C1 => IR_IN(27), C2 => n13, A => n15, B => n12, ZN
                           => cw_1_port);
   U14 : NAND3_X1 port map( A1 => n16, A2 => n4, A3 => n17, ZN => cw_17_port);
   U15 : NAND4_X1 port map( A1 => n8, A2 => n9, A3 => n18, A4 => n19, ZN => n16
                           );
   U16 : OR2_X1 port map( A1 => cw_6_port, A2 => n20, ZN => cw_14_port);
   U17 : NOR4_X1 port map( A1 => n21, A2 => n22, A3 => n9, A4 => n18, ZN => 
                           cw_6_port);
   U18 : INV_X1 port map( A => IR_IN(29), ZN => n22);
   U19 : OAI211_X1 port map( C1 => IR_IN(30), C2 => n4, A => n15, B => n17, ZN 
                           => cw_13_port);
   U20 : AND3_X1 port map( A1 => n10, A2 => n7, A3 => n12, ZN => n17);
   U21 : NOR3_X1 port map( A1 => n23, A2 => n24, A3 => n25, ZN => n12);
   U22 : NAND4_X1 port map( A1 => n26, A2 => n27, A3 => n28, A4 => n13, ZN => 
                           cw_12_port);
   U23 : AND2_X1 port map( A1 => n11, A2 => n10, ZN => n28);
   U24 : NAND4_X1 port map( A1 => IR_IN(30), A2 => IR_IN(28), A3 => IR_IN(29), 
                           A4 => n18, ZN => n26);
   U25 : OAI211_X1 port map( C1 => IR_IN(31), C2 => n29, A => n30, B => n31, ZN
                           => aluOpcode_i_3_port);
   U26 : NAND3_X1 port map( A1 => IR_IN(3), A2 => IR_IN(0), A3 => n32, ZN => 
                           n30);
   U27 : NOR3_X1 port map( A1 => n33, A2 => IR_IN(2), A3 => IR_IN(1), ZN => n32
                           );
   U28 : AOI21_X1 port map( B1 => n25, B2 => n19, A => n23, ZN => n29);
   U29 : INV_X1 port map( A => n27, ZN => n25);
   U30 : NAND3_X1 port map( A1 => IR_IN(29), A2 => n18, A3 => n3, ZN => n27);
   U31 : OAI221_X1 port map( B1 => n35, B2 => n36, C1 => n37, C2 => n15, A => 
                           n38, ZN => aluOpcode_i_2_port);
   U32 : AOI211_X1 port map( C1 => n39, C2 => IR_IN(1), A => n40, B => n41, ZN 
                           => n38);
   U33 : NOR3_X1 port map( A1 => n42, A2 => n18, A3 => n19, ZN => n40);
   U34 : NOR2_X1 port map( A1 => n43, A2 => n44, ZN => n39);
   U35 : INV_X1 port map( A => n45, ZN => n36);
   U36 : NAND4_X1 port map( A1 => n46, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           aluOpcode_i_1_port);
   U37 : AOI221_X1 port map( B1 => n45, B2 => n35, C1 => n24, C2 => n14, A => 
                           n50, ZN => n49);
   U38 : MUX2_X1 port map( A => n51, B => n52, S => IR_IN(1), Z => n50);
   U39 : NOR3_X1 port map( A1 => n44, A2 => IR_IN(2), A3 => n33, ZN => n52);
   U40 : INV_X1 port map( A => n53, ZN => n44);
   U41 : INV_X1 port map( A => n42, ZN => n24);
   U42 : INV_X1 port map( A => IR_IN(0), ZN => n35);
   U43 : OR3_X1 port map( A1 => n8, A2 => IR_IN(26), A3 => n4, ZN => n48);
   U44 : NAND4_X1 port map( A1 => n46, A2 => n11, A3 => n54, A4 => n55, ZN => 
                           aluOpcode_i_0_port);
   U45 : AOI221_X1 port map( B1 => n41, B2 => IR_IN(0), C1 => n51, C2 => 
                           IR_IN(1), A => n56, ZN => n55);
   U46 : OAI22_X1 port map( A1 => n14, A2 => n42, B1 => IR_IN(30), B2 => n10, 
                           ZN => n56);
   U47 : NAND3_X1 port map( A1 => IR_IN(26), A2 => n14, A3 => IR_IN(31), ZN => 
                           n10);
   U48 : NAND3_X1 port map( A1 => n37, A2 => n21, A3 => IR_IN(29), ZN => n42);
   U49 : INV_X1 port map( A => n31, ZN => n51);
   U50 : NAND4_X1 port map( A1 => n20, A2 => n57, A3 => IR_IN(2), A4 => n58, ZN
                           => n31);
   U51 : NOR3_X1 port map( A1 => IR_IN(0), A2 => IR_IN(5), A3 => IR_IN(3), ZN 
                           => n58);
   U52 : INV_X1 port map( A => n47, ZN => n41);
   U53 : NAND2_X1 port map( A1 => n45, A2 => IR_IN(3), ZN => n47);
   U54 : NOR2_X1 port map( A1 => n43, A2 => IR_IN(1), ZN => n45);
   U55 : AOI21_X1 port map( B1 => n53, B2 => n59, A => n60, ZN => n54);
   U56 : AND3_X1 port map( A1 => n23, A2 => n21, A3 => IR_IN(27), ZN => n60);
   U57 : NOR4_X1 port map( A1 => n61, A2 => n19, A3 => IR_IN(26), A4 => 
                           IR_IN(29), ZN => n23);
   U58 : OAI21_X1 port map( B1 => IR_IN(1), B2 => n33, A => n43, ZN => n59);
   U59 : NAND2_X1 port map( A1 => n62, A2 => IR_IN(2), ZN => n43);
   U60 : INV_X1 port map( A => n33, ZN => n62);
   U61 : NAND3_X1 port map( A1 => n20, A2 => n57, A3 => IR_IN(5), ZN => n33);
   U62 : NOR4_X1 port map( A1 => IR_IN(6), A2 => IR_IN(4), A3 => IR_IN(10), A4 
                           => n63, ZN => n57);
   U63 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN =>
                           n63);
   U64 : NOR3_X1 port map( A1 => IR_IN(27), A2 => IR_IN(29), A3 => n13, ZN => 
                           n20);
   U65 : NAND3_X1 port map( A1 => n19, A2 => n21, A3 => n37, ZN => n13);
   U66 : NOR2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(26), ZN => n37);
   U67 : INV_X1 port map( A => IR_IN(28), ZN => n19);
   U68 : NOR2_X1 port map( A1 => IR_IN(0), A2 => IR_IN(3), ZN => n53);
   U69 : AOI21_X1 port map( B1 => n8, B2 => n64, A => n66, ZN => n11);
   U70 : INV_X1 port map( A => n7, ZN => n66);
   U71 : NAND3_X1 port map( A1 => n8, A2 => n21, A3 => n14, ZN => n7);
   U72 : NOR2_X1 port map( A1 => n18, A2 => IR_IN(28), ZN => n14);
   U73 : NOR2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), ZN => n8);
   U74 : NAND2_X1 port map( A1 => n65, A2 => n3, ZN => n46);
   U75 : NOR2_X1 port map( A1 => n61, A2 => n9, ZN => n3);
   U76 : INV_X1 port map( A => IR_IN(26), ZN => n9);
   U77 : INV_X1 port map( A => IR_IN(30), ZN => n61);
   U78 : INV_X1 port map( A => n15, ZN => n65);
   U79 : NAND2_X1 port map( A1 => n64, A2 => IR_IN(29), ZN => n15);
   U80 : INV_X1 port map( A => n4, ZN => n64);
   U81 : NAND3_X1 port map( A1 => n18, A2 => n21, A3 => IR_IN(28), ZN => n4);
   U82 : INV_X1 port map( A => IR_IN(31), ZN => n21);
   U83 : INV_X1 port map( A => IR_IN(27), ZN => n18);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 is

   port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
         EQ_COND, IS_JUMP : in std_logic;  ALU_OPCODE : in std_logic_vector (0 
         to 3);  JUMP_EN, PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE : in std_logic
         ;  D_ADDR : out std_logic_vector (5 downto 0);  D_DATA_IN : out 
         std_logic_vector (31 downto 0);  D_DATA_OUT, PC_IN : in 
         std_logic_vector (31 downto 0);  PC_BUS : out std_logic_vector (31 
         downto 0));

end DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64;

architecture SYN_STRUCTURE of 
   DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component ALU_N32
      port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26
      port( NOT_EXT_IMM : in std_logic_vector (25 downto 0);  SIGNED_IMM, 
            IS_JUMP : in std_logic;  EXT_IMM : out std_logic_vector (31 downto 
            0));
   end component;
   
   component REGISTER_FILE_NBIT32_NREG32
      port( CLK, RST, EN, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component ADDER_N32
      port( CURR_ADDR : in std_logic_vector (31 downto 0);  NEXT_ADDR : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT5_1
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT5_0
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component MUX21
      port( A, B, SEL : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component BRANCHING_UNIT_N32
      port( CLK, RST : in std_logic;  Reg_A : in std_logic_vector (31 downto 0)
            ;  EQ_cond, IS_JUMP : in std_logic;  branch_taken : out std_logic);
   end component;
   
   component REG_GENERIC_NBIT32_1
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_2
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_3
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT5_1
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 
            downto 0);  DATA_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component REG_GENERIC_NBIT5_2
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 
            downto 0);  DATA_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component REG_GENERIC_NBIT5_0
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (4 
            downto 0);  DATA_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component REG_GENERIC_NBIT26
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (25 
            downto 0);  DATA_OUT : out std_logic_vector (25 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_4
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_5
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_6
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_7
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_8
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, D_ADDR_5_port, D_ADDR_4_port, 
      D_ADDR_3_port, D_ADDR_2_port, D_ADDR_1_port, D_ADDR_0_port, 
      PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, current_PC_31_port, 
      current_PC_30_port, current_PC_29_port, current_PC_28_port, 
      current_PC_27_port, current_PC_26_port, current_PC_25_port, 
      current_PC_24_port, current_PC_23_port, current_PC_22_port, 
      current_PC_21_port, current_PC_20_port, current_PC_19_port, 
      current_PC_18_port, current_PC_17_port, current_PC_16_port, 
      current_PC_15_port, current_PC_14_port, current_PC_13_port, 
      current_PC_12_port, current_PC_11_port, current_PC_10_port, 
      current_PC_9_port, current_PC_8_port, current_PC_7_port, 
      current_PC_6_port, current_PC_5_port, current_PC_4_port, 
      current_PC_3_port, current_PC_2_port, current_PC_1_port, 
      current_PC_0_port, current_PC1_31_port, current_PC1_30_port, 
      current_PC1_29_port, current_PC1_28_port, current_PC1_27_port, 
      current_PC1_26_port, current_PC1_25_port, current_PC1_24_port, 
      current_PC1_23_port, current_PC1_22_port, current_PC1_21_port, 
      current_PC1_20_port, current_PC1_19_port, current_PC1_18_port, 
      current_PC1_17_port, current_PC1_16_port, current_PC1_15_port, 
      current_PC1_14_port, current_PC1_13_port, current_PC1_12_port, 
      current_PC1_11_port, current_PC1_10_port, current_PC1_9_port, 
      current_PC1_8_port, current_PC1_7_port, current_PC1_6_port, 
      current_PC1_5_port, current_PC1_4_port, current_PC1_3_port, 
      current_PC1_2_port, current_PC1_1_port, current_PC1_0_port, 
      current_PC2_31_port, current_PC2_30_port, current_PC2_29_port, 
      current_PC2_28_port, current_PC2_27_port, current_PC2_26_port, 
      current_PC2_25_port, current_PC2_24_port, current_PC2_23_port, 
      current_PC2_22_port, current_PC2_21_port, current_PC2_20_port, 
      current_PC2_19_port, current_PC2_18_port, current_PC2_17_port, 
      current_PC2_16_port, current_PC2_15_port, current_PC2_14_port, 
      current_PC2_13_port, current_PC2_12_port, current_PC2_11_port, 
      current_PC2_10_port, current_PC2_9_port, current_PC2_8_port, 
      current_PC2_7_port, current_PC2_6_port, current_PC2_5_port, 
      current_PC2_4_port, current_PC2_3_port, current_PC2_2_port, 
      current_PC2_1_port, current_PC2_0_port, current_PC3_31_port, 
      current_PC3_30_port, current_PC3_29_port, current_PC3_28_port, 
      current_PC3_27_port, current_PC3_26_port, current_PC3_25_port, 
      current_PC3_24_port, current_PC3_23_port, current_PC3_22_port, 
      current_PC3_21_port, current_PC3_20_port, current_PC3_19_port, 
      current_PC3_18_port, current_PC3_17_port, current_PC3_16_port, 
      current_PC3_15_port, current_PC3_14_port, current_PC3_13_port, 
      current_PC3_12_port, current_PC3_11_port, current_PC3_10_port, 
      current_PC3_9_port, current_PC3_8_port, current_PC3_7_port, 
      current_PC3_6_port, current_PC3_5_port, current_PC3_4_port, 
      current_PC3_3_port, current_PC3_2_port, current_PC3_1_port, 
      current_PC3_0_port, next_NPC_31_port, next_NPC_30_port, next_NPC_29_port,
      next_NPC_28_port, next_NPC_27_port, next_NPC_26_port, next_NPC_25_port, 
      next_NPC_24_port, next_NPC_23_port, next_NPC_22_port, next_NPC_21_port, 
      next_NPC_20_port, next_NPC_19_port, next_NPC_18_port, next_NPC_17_port, 
      next_NPC_16_port, next_NPC_15_port, next_NPC_14_port, next_NPC_13_port, 
      next_NPC_12_port, next_NPC_11_port, next_NPC_10_port, next_NPC_9_port, 
      next_NPC_8_port, next_NPC_7_port, next_NPC_6_port, next_NPC_5_port, 
      next_NPC_4_port, next_NPC_3_port, next_NPC_2_port, next_NPC_1_port, 
      next_NPC_0_port, current_NPC_31_port, current_NPC_30_port, 
      current_NPC_29_port, current_NPC_28_port, current_NPC_27_port, 
      current_NPC_26_port, current_NPC_25_port, current_NPC_24_port, 
      current_NPC_23_port, current_NPC_22_port, current_NPC_21_port, 
      current_NPC_20_port, current_NPC_19_port, current_NPC_18_port, 
      current_NPC_17_port, current_NPC_16_port, current_NPC_15_port, 
      current_NPC_14_port, current_NPC_13_port, current_NPC_12_port, 
      current_NPC_11_port, current_NPC_10_port, current_NPC_9_port, 
      current_NPC_8_port, current_NPC_7_port, current_NPC_6_port, 
      current_NPC_5_port, current_NPC_4_port, current_NPC_3_port, 
      current_NPC_2_port, current_NPC_1_port, current_NPC_0_port, 
      current_IW_25_port, current_IW_24_port, current_IW_23_port, 
      current_IW_22_port, current_IW_21_port, current_IW_20_port, 
      current_IW_19_port, current_IW_18_port, current_IW_17_port, 
      current_IW_16_port, current_IW_15_port, current_IW_14_port, 
      current_IW_13_port, current_IW_12_port, current_IW_11_port, 
      current_IW_10_port, current_IW_9_port, current_IW_8_port, 
      current_IW_7_port, current_IW_6_port, current_IW_5_port, 
      current_IW_4_port, current_IW_3_port, current_IW_2_port, 
      current_IW_1_port, current_IW_0_port, IMM_IN_25_port, IMM_IN_24_port, 
      IMM_IN_23_port, IMM_IN_22_port, IMM_IN_21_port, IMM_IN_20_port, 
      IMM_IN_19_port, IMM_IN_18_port, IMM_IN_17_port, IMM_IN_16_port, 
      IMM_IN_15_port, IMM_IN_14_port, IMM_IN_13_port, IMM_IN_12_port, 
      IMM_IN_11_port, IMM_IN_10_port, IMM_IN_9_port, IMM_IN_8_port, 
      IMM_IN_7_port, IMM_IN_6_port, IMM_IN_5_port, IMM_IN_4_port, IMM_IN_3_port
      , IMM_IN_2_port, IMM_IN_1_port, IMM_IN_0_port, WB1_IN_4_port, 
      WB1_IN_3_port, WB1_IN_2_port, WB1_IN_1_port, WB1_IN_0_port, WB2_IN_4_port
      , WB2_IN_3_port, WB2_IN_2_port, WB2_IN_1_port, WB2_IN_0_port, 
      WB2_OUT_4_port, WB2_OUT_3_port, WB2_OUT_2_port, WB2_OUT_1_port, 
      WB2_OUT_0_port, WB3_OUT_4_port, WB3_OUT_3_port, WB3_OUT_2_port, 
      WB3_OUT_1_port, WB3_OUT_0_port, next_ALU_OUT_31_port, 
      next_ALU_OUT_30_port, next_ALU_OUT_29_port, next_ALU_OUT_28_port, 
      next_ALU_OUT_27_port, next_ALU_OUT_26_port, next_ALU_OUT_25_port, 
      next_ALU_OUT_24_port, next_ALU_OUT_23_port, next_ALU_OUT_22_port, 
      next_ALU_OUT_21_port, next_ALU_OUT_20_port, next_ALU_OUT_19_port, 
      next_ALU_OUT_18_port, next_ALU_OUT_17_port, next_ALU_OUT_16_port, 
      next_ALU_OUT_15_port, next_ALU_OUT_14_port, next_ALU_OUT_13_port, 
      next_ALU_OUT_12_port, next_ALU_OUT_11_port, next_ALU_OUT_10_port, 
      next_ALU_OUT_9_port, next_ALU_OUT_8_port, next_ALU_OUT_7_port, 
      next_ALU_OUT_6_port, next_ALU_OUT_5_port, next_ALU_OUT_4_port, 
      next_ALU_OUT_3_port, next_ALU_OUT_2_port, next_ALU_OUT_1_port, 
      next_ALU_OUT_0_port, current_ALU_OUT_31_port, current_ALU_OUT_30_port, 
      current_ALU_OUT_29_port, current_ALU_OUT_28_port, current_ALU_OUT_27_port
      , current_ALU_OUT_26_port, current_ALU_OUT_25_port, 
      current_ALU_OUT_24_port, current_ALU_OUT_23_port, current_ALU_OUT_22_port
      , current_ALU_OUT_21_port, current_ALU_OUT_20_port, 
      current_ALU_OUT_19_port, current_ALU_OUT_18_port, current_ALU_OUT_17_port
      , current_ALU_OUT_16_port, current_ALU_OUT_15_port, 
      current_ALU_OUT_14_port, current_ALU_OUT_13_port, current_ALU_OUT_12_port
      , current_ALU_OUT_11_port, current_ALU_OUT_10_port, 
      current_ALU_OUT_9_port, current_ALU_OUT_8_port, current_ALU_OUT_7_port, 
      current_ALU_OUT_6_port, B_OUT_31_port, B_OUT_30_port, B_OUT_29_port, 
      B_OUT_28_port, B_OUT_27_port, B_OUT_26_port, B_OUT_25_port, B_OUT_24_port
      , B_OUT_23_port, B_OUT_22_port, B_OUT_21_port, B_OUT_20_port, 
      B_OUT_19_port, B_OUT_18_port, B_OUT_17_port, B_OUT_16_port, B_OUT_15_port
      , B_OUT_14_port, B_OUT_13_port, B_OUT_12_port, B_OUT_11_port, 
      B_OUT_10_port, B_OUT_9_port, B_OUT_8_port, B_OUT_7_port, B_OUT_6_port, 
      B_OUT_5_port, B_OUT_4_port, B_OUT_3_port, B_OUT_2_port, B_OUT_1_port, 
      B_OUT_0_port, current_ALU_OUT2_31_port, current_ALU_OUT2_30_port, 
      current_ALU_OUT2_29_port, current_ALU_OUT2_28_port, 
      current_ALU_OUT2_27_port, current_ALU_OUT2_26_port, 
      current_ALU_OUT2_25_port, current_ALU_OUT2_24_port, 
      current_ALU_OUT2_23_port, current_ALU_OUT2_22_port, 
      current_ALU_OUT2_21_port, current_ALU_OUT2_20_port, 
      current_ALU_OUT2_19_port, current_ALU_OUT2_18_port, 
      current_ALU_OUT2_17_port, current_ALU_OUT2_16_port, 
      current_ALU_OUT2_15_port, current_ALU_OUT2_14_port, 
      current_ALU_OUT2_13_port, current_ALU_OUT2_12_port, 
      current_ALU_OUT2_11_port, current_ALU_OUT2_10_port, 
      current_ALU_OUT2_9_port, current_ALU_OUT2_8_port, current_ALU_OUT2_7_port
      , current_ALU_OUT2_6_port, current_ALU_OUT2_5_port, 
      current_ALU_OUT2_4_port, current_ALU_OUT2_3_port, current_ALU_OUT2_2_port
      , current_ALU_OUT2_1_port, current_ALU_OUT2_0_port, A_OUT_31_port, 
      A_OUT_30_port, A_OUT_29_port, A_OUT_28_port, A_OUT_27_port, A_OUT_26_port
      , A_OUT_25_port, A_OUT_24_port, A_OUT_23_port, A_OUT_22_port, 
      A_OUT_21_port, A_OUT_20_port, A_OUT_19_port, A_OUT_18_port, A_OUT_17_port
      , A_OUT_16_port, A_OUT_15_port, A_OUT_14_port, A_OUT_13_port, 
      A_OUT_12_port, A_OUT_11_port, A_OUT_10_port, A_OUT_9_port, A_OUT_8_port, 
      A_OUT_7_port, A_OUT_6_port, A_OUT_5_port, A_OUT_4_port, A_OUT_3_port, 
      A_OUT_2_port, A_OUT_1_port, A_OUT_0_port, branch_taken, PC_MUX_SEL, 
      ALU_OP1_31_port, ALU_OP1_30_port, ALU_OP1_29_port, ALU_OP1_28_port, 
      ALU_OP1_27_port, ALU_OP1_26_port, ALU_OP1_25_port, ALU_OP1_24_port, 
      ALU_OP1_23_port, ALU_OP1_22_port, ALU_OP1_21_port, ALU_OP1_20_port, 
      ALU_OP1_19_port, ALU_OP1_18_port, ALU_OP1_17_port, ALU_OP1_16_port, 
      ALU_OP1_15_port, ALU_OP1_14_port, ALU_OP1_13_port, ALU_OP1_12_port, 
      ALU_OP1_11_port, ALU_OP1_10_port, ALU_OP1_9_port, ALU_OP1_8_port, 
      ALU_OP1_7_port, ALU_OP1_6_port, ALU_OP1_5_port, ALU_OP1_4_port, 
      ALU_OP1_3_port, ALU_OP1_2_port, ALU_OP1_1_port, ALU_OP1_0_port, 
      IMM_OUT_31_port, IMM_OUT_30_port, IMM_OUT_29_port, IMM_OUT_28_port, 
      IMM_OUT_27_port, IMM_OUT_26_port, IMM_OUT_25_port, IMM_OUT_24_port, 
      IMM_OUT_23_port, IMM_OUT_22_port, IMM_OUT_21_port, IMM_OUT_20_port, 
      IMM_OUT_19_port, IMM_OUT_18_port, IMM_OUT_17_port, IMM_OUT_16_port, 
      IMM_OUT_15_port, IMM_OUT_14_port, IMM_OUT_13_port, IMM_OUT_12_port, 
      IMM_OUT_11_port, IMM_OUT_10_port, IMM_OUT_9_port, IMM_OUT_8_port, 
      IMM_OUT_7_port, IMM_OUT_6_port, IMM_OUT_5_port, IMM_OUT_4_port, 
      IMM_OUT_3_port, IMM_OUT_2_port, IMM_OUT_1_port, IMM_OUT_0_port, 
      ALU_OP2_31_port, ALU_OP2_30_port, ALU_OP2_29_port, ALU_OP2_28_port, 
      ALU_OP2_27_port, ALU_OP2_26_port, ALU_OP2_25_port, ALU_OP2_24_port, 
      ALU_OP2_23_port, ALU_OP2_22_port, ALU_OP2_21_port, ALU_OP2_20_port, 
      ALU_OP2_19_port, ALU_OP2_18_port, ALU_OP2_17_port, ALU_OP2_16_port, 
      ALU_OP2_15_port, ALU_OP2_14_port, ALU_OP2_13_port, ALU_OP2_12_port, 
      ALU_OP2_11_port, ALU_OP2_10_port, ALU_OP2_9_port, ALU_OP2_8_port, 
      ALU_OP2_7_port, ALU_OP2_6_port, ALU_OP2_5_port, ALU_OP2_4_port, 
      ALU_OP2_3_port, ALU_OP2_2_port, ALU_OP2_1_port, ALU_OP2_0_port, 
      OUT_MUX_DATA_31_port, OUT_MUX_DATA_30_port, OUT_MUX_DATA_29_port, 
      OUT_MUX_DATA_28_port, OUT_MUX_DATA_27_port, OUT_MUX_DATA_26_port, 
      OUT_MUX_DATA_25_port, OUT_MUX_DATA_24_port, OUT_MUX_DATA_23_port, 
      OUT_MUX_DATA_22_port, OUT_MUX_DATA_21_port, OUT_MUX_DATA_20_port, 
      OUT_MUX_DATA_19_port, OUT_MUX_DATA_18_port, OUT_MUX_DATA_17_port, 
      OUT_MUX_DATA_16_port, OUT_MUX_DATA_15_port, OUT_MUX_DATA_14_port, 
      OUT_MUX_DATA_13_port, OUT_MUX_DATA_12_port, OUT_MUX_DATA_11_port, 
      OUT_MUX_DATA_10_port, OUT_MUX_DATA_9_port, OUT_MUX_DATA_8_port, 
      OUT_MUX_DATA_7_port, OUT_MUX_DATA_6_port, OUT_MUX_DATA_5_port, 
      OUT_MUX_DATA_4_port, OUT_MUX_DATA_3_port, OUT_MUX_DATA_2_port, 
      OUT_MUX_DATA_1_port, OUT_MUX_DATA_0_port, WB_DATA_31_port, 
      WB_DATA_30_port, WB_DATA_29_port, WB_DATA_28_port, WB_DATA_27_port, 
      WB_DATA_26_port, WB_DATA_25_port, WB_DATA_24_port, WB_DATA_23_port, 
      WB_DATA_22_port, WB_DATA_21_port, WB_DATA_20_port, WB_DATA_19_port, 
      WB_DATA_18_port, WB_DATA_17_port, WB_DATA_16_port, WB_DATA_15_port, 
      WB_DATA_14_port, WB_DATA_13_port, WB_DATA_12_port, WB_DATA_11_port, 
      WB_DATA_10_port, WB_DATA_9_port, WB_DATA_8_port, WB_DATA_7_port, 
      WB_DATA_6_port, WB_DATA_5_port, WB_DATA_4_port, WB_DATA_3_port, 
      WB_DATA_2_port, WB_DATA_1_port, WB_DATA_0_port, WB_ADDR_4_port, 
      WB_ADDR_3_port, WB_ADDR_2_port, WB_ADDR_1_port, WB_ADDR_0_port, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612 : std_logic;

begin
   D_ADDR <= ( D_ADDR_5_port, D_ADDR_4_port, D_ADDR_3_port, D_ADDR_2_port, 
      D_ADDR_1_port, D_ADDR_0_port );
   PC_BUS <= ( PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   PC_REG : REG_GENERIC_NBIT32_8 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => PC_IN(31), DATA_IN(30) 
                           => PC_IN(30), DATA_IN(29) => PC_IN(29), DATA_IN(28) 
                           => PC_IN(28), DATA_IN(27) => PC_IN(27), DATA_IN(26) 
                           => PC_IN(26), DATA_IN(25) => PC_IN(25), DATA_IN(24) 
                           => PC_IN(24), DATA_IN(23) => PC_IN(23), DATA_IN(22) 
                           => PC_IN(22), DATA_IN(21) => PC_IN(21), DATA_IN(20) 
                           => PC_IN(20), DATA_IN(19) => PC_IN(19), DATA_IN(18) 
                           => PC_IN(18), DATA_IN(17) => PC_IN(17), DATA_IN(16) 
                           => PC_IN(16), DATA_IN(15) => PC_IN(15), DATA_IN(14) 
                           => PC_IN(14), DATA_IN(13) => PC_IN(13), DATA_IN(12) 
                           => PC_IN(12), DATA_IN(11) => PC_IN(11), DATA_IN(10) 
                           => PC_IN(10), DATA_IN(9) => PC_IN(9), DATA_IN(8) => 
                           PC_IN(8), DATA_IN(7) => PC_IN(7), DATA_IN(6) => 
                           PC_IN(6), DATA_IN(5) => PC_IN(5), DATA_IN(4) => 
                           PC_IN(4), DATA_IN(3) => PC_IN(3), DATA_IN(2) => 
                           PC_IN(2), DATA_IN(1) => PC_IN(1), DATA_IN(0) => 
                           PC_IN(0), DATA_OUT(31) => current_PC1_31_port, 
                           DATA_OUT(30) => current_PC1_30_port, DATA_OUT(29) =>
                           current_PC1_29_port, DATA_OUT(28) => 
                           current_PC1_28_port, DATA_OUT(27) => 
                           current_PC1_27_port, DATA_OUT(26) => 
                           current_PC1_26_port, DATA_OUT(25) => 
                           current_PC1_25_port, DATA_OUT(24) => 
                           current_PC1_24_port, DATA_OUT(23) => 
                           current_PC1_23_port, DATA_OUT(22) => 
                           current_PC1_22_port, DATA_OUT(21) => 
                           current_PC1_21_port, DATA_OUT(20) => 
                           current_PC1_20_port, DATA_OUT(19) => 
                           current_PC1_19_port, DATA_OUT(18) => 
                           current_PC1_18_port, DATA_OUT(17) => 
                           current_PC1_17_port, DATA_OUT(16) => 
                           current_PC1_16_port, DATA_OUT(15) => 
                           current_PC1_15_port, DATA_OUT(14) => 
                           current_PC1_14_port, DATA_OUT(13) => 
                           current_PC1_13_port, DATA_OUT(12) => 
                           current_PC1_12_port, DATA_OUT(11) => 
                           current_PC1_11_port, DATA_OUT(10) => 
                           current_PC1_10_port, DATA_OUT(9) => 
                           current_PC1_9_port, DATA_OUT(8) => 
                           current_PC1_8_port, DATA_OUT(7) => 
                           current_PC1_7_port, DATA_OUT(6) => 
                           current_PC1_6_port, DATA_OUT(5) => 
                           current_PC1_5_port, DATA_OUT(4) => 
                           current_PC1_4_port, DATA_OUT(3) => 
                           current_PC1_3_port, DATA_OUT(2) => 
                           current_PC1_2_port, DATA_OUT(1) => 
                           current_PC1_1_port, DATA_OUT(0) => 
                           current_PC1_0_port);
   PC2_REG : REG_GENERIC_NBIT32_7 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => current_PC1_31_port, 
                           DATA_IN(30) => current_PC1_30_port, DATA_IN(29) => 
                           current_PC1_29_port, DATA_IN(28) => 
                           current_PC1_28_port, DATA_IN(27) => 
                           current_PC1_27_port, DATA_IN(26) => 
                           current_PC1_26_port, DATA_IN(25) => 
                           current_PC1_25_port, DATA_IN(24) => 
                           current_PC1_24_port, DATA_IN(23) => 
                           current_PC1_23_port, DATA_IN(22) => 
                           current_PC1_22_port, DATA_IN(21) => 
                           current_PC1_21_port, DATA_IN(20) => 
                           current_PC1_20_port, DATA_IN(19) => 
                           current_PC1_19_port, DATA_IN(18) => 
                           current_PC1_18_port, DATA_IN(17) => 
                           current_PC1_17_port, DATA_IN(16) => 
                           current_PC1_16_port, DATA_IN(15) => 
                           current_PC1_15_port, DATA_IN(14) => 
                           current_PC1_14_port, DATA_IN(13) => 
                           current_PC1_13_port, DATA_IN(12) => 
                           current_PC1_12_port, DATA_IN(11) => 
                           current_PC1_11_port, DATA_IN(10) => 
                           current_PC1_10_port, DATA_IN(9) => 
                           current_PC1_9_port, DATA_IN(8) => current_PC1_8_port
                           , DATA_IN(7) => current_PC1_7_port, DATA_IN(6) => 
                           current_PC1_6_port, DATA_IN(5) => current_PC1_5_port
                           , DATA_IN(4) => current_PC1_4_port, DATA_IN(3) => 
                           current_PC1_3_port, DATA_IN(2) => current_PC1_2_port
                           , DATA_IN(1) => current_PC1_1_port, DATA_IN(0) => 
                           current_PC1_0_port, DATA_OUT(31) => 
                           current_PC2_31_port, DATA_OUT(30) => 
                           current_PC2_30_port, DATA_OUT(29) => 
                           current_PC2_29_port, DATA_OUT(28) => 
                           current_PC2_28_port, DATA_OUT(27) => 
                           current_PC2_27_port, DATA_OUT(26) => 
                           current_PC2_26_port, DATA_OUT(25) => 
                           current_PC2_25_port, DATA_OUT(24) => 
                           current_PC2_24_port, DATA_OUT(23) => 
                           current_PC2_23_port, DATA_OUT(22) => 
                           current_PC2_22_port, DATA_OUT(21) => 
                           current_PC2_21_port, DATA_OUT(20) => 
                           current_PC2_20_port, DATA_OUT(19) => 
                           current_PC2_19_port, DATA_OUT(18) => 
                           current_PC2_18_port, DATA_OUT(17) => 
                           current_PC2_17_port, DATA_OUT(16) => 
                           current_PC2_16_port, DATA_OUT(15) => 
                           current_PC2_15_port, DATA_OUT(14) => 
                           current_PC2_14_port, DATA_OUT(13) => 
                           current_PC2_13_port, DATA_OUT(12) => 
                           current_PC2_12_port, DATA_OUT(11) => 
                           current_PC2_11_port, DATA_OUT(10) => 
                           current_PC2_10_port, DATA_OUT(9) => 
                           current_PC2_9_port, DATA_OUT(8) => 
                           current_PC2_8_port, DATA_OUT(7) => 
                           current_PC2_7_port, DATA_OUT(6) => 
                           current_PC2_6_port, DATA_OUT(5) => 
                           current_PC2_5_port, DATA_OUT(4) => 
                           current_PC2_4_port, DATA_OUT(3) => 
                           current_PC2_3_port, DATA_OUT(2) => 
                           current_PC2_2_port, DATA_OUT(1) => 
                           current_PC2_1_port, DATA_OUT(0) => 
                           current_PC2_0_port);
   PC3_REG : REG_GENERIC_NBIT32_6 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => current_PC2_31_port, 
                           DATA_IN(30) => current_PC2_30_port, DATA_IN(29) => 
                           current_PC2_29_port, DATA_IN(28) => 
                           current_PC2_28_port, DATA_IN(27) => 
                           current_PC2_27_port, DATA_IN(26) => 
                           current_PC2_26_port, DATA_IN(25) => 
                           current_PC2_25_port, DATA_IN(24) => 
                           current_PC2_24_port, DATA_IN(23) => 
                           current_PC2_23_port, DATA_IN(22) => 
                           current_PC2_22_port, DATA_IN(21) => 
                           current_PC2_21_port, DATA_IN(20) => 
                           current_PC2_20_port, DATA_IN(19) => 
                           current_PC2_19_port, DATA_IN(18) => 
                           current_PC2_18_port, DATA_IN(17) => 
                           current_PC2_17_port, DATA_IN(16) => 
                           current_PC2_16_port, DATA_IN(15) => 
                           current_PC2_15_port, DATA_IN(14) => 
                           current_PC2_14_port, DATA_IN(13) => 
                           current_PC2_13_port, DATA_IN(12) => 
                           current_PC2_12_port, DATA_IN(11) => 
                           current_PC2_11_port, DATA_IN(10) => 
                           current_PC2_10_port, DATA_IN(9) => 
                           current_PC2_9_port, DATA_IN(8) => current_PC2_8_port
                           , DATA_IN(7) => current_PC2_7_port, DATA_IN(6) => 
                           current_PC2_6_port, DATA_IN(5) => current_PC2_5_port
                           , DATA_IN(4) => current_PC2_4_port, DATA_IN(3) => 
                           current_PC2_3_port, DATA_IN(2) => current_PC2_2_port
                           , DATA_IN(1) => current_PC2_1_port, DATA_IN(0) => 
                           current_PC2_0_port, DATA_OUT(31) => 
                           current_PC3_31_port, DATA_OUT(30) => 
                           current_PC3_30_port, DATA_OUT(29) => 
                           current_PC3_29_port, DATA_OUT(28) => 
                           current_PC3_28_port, DATA_OUT(27) => 
                           current_PC3_27_port, DATA_OUT(26) => 
                           current_PC3_26_port, DATA_OUT(25) => 
                           current_PC3_25_port, DATA_OUT(24) => 
                           current_PC3_24_port, DATA_OUT(23) => 
                           current_PC3_23_port, DATA_OUT(22) => 
                           current_PC3_22_port, DATA_OUT(21) => 
                           current_PC3_21_port, DATA_OUT(20) => 
                           current_PC3_20_port, DATA_OUT(19) => 
                           current_PC3_19_port, DATA_OUT(18) => 
                           current_PC3_18_port, DATA_OUT(17) => 
                           current_PC3_17_port, DATA_OUT(16) => 
                           current_PC3_16_port, DATA_OUT(15) => 
                           current_PC3_15_port, DATA_OUT(14) => 
                           current_PC3_14_port, DATA_OUT(13) => 
                           current_PC3_13_port, DATA_OUT(12) => 
                           current_PC3_12_port, DATA_OUT(11) => 
                           current_PC3_11_port, DATA_OUT(10) => 
                           current_PC3_10_port, DATA_OUT(9) => 
                           current_PC3_9_port, DATA_OUT(8) => 
                           current_PC3_8_port, DATA_OUT(7) => 
                           current_PC3_7_port, DATA_OUT(6) => 
                           current_PC3_6_port, DATA_OUT(5) => 
                           current_PC3_5_port, DATA_OUT(4) => 
                           current_PC3_4_port, DATA_OUT(3) => 
                           current_PC3_3_port, DATA_OUT(2) => 
                           current_PC3_2_port, DATA_OUT(1) => 
                           current_PC3_1_port, DATA_OUT(0) => 
                           current_PC3_0_port);
   NPC_REG : REG_GENERIC_NBIT32_5 port map( CLK => CLK, RST => RST, EN => 
                           NPC_LATCH_EN, DATA_IN(31) => next_NPC_31_port, 
                           DATA_IN(30) => next_NPC_30_port, DATA_IN(29) => 
                           next_NPC_29_port, DATA_IN(28) => next_NPC_28_port, 
                           DATA_IN(27) => next_NPC_27_port, DATA_IN(26) => 
                           next_NPC_26_port, DATA_IN(25) => next_NPC_25_port, 
                           DATA_IN(24) => next_NPC_24_port, DATA_IN(23) => 
                           next_NPC_23_port, DATA_IN(22) => next_NPC_22_port, 
                           DATA_IN(21) => next_NPC_21_port, DATA_IN(20) => 
                           next_NPC_20_port, DATA_IN(19) => next_NPC_19_port, 
                           DATA_IN(18) => next_NPC_18_port, DATA_IN(17) => 
                           next_NPC_17_port, DATA_IN(16) => next_NPC_16_port, 
                           DATA_IN(15) => next_NPC_15_port, DATA_IN(14) => 
                           next_NPC_14_port, DATA_IN(13) => next_NPC_13_port, 
                           DATA_IN(12) => next_NPC_12_port, DATA_IN(11) => 
                           next_NPC_11_port, DATA_IN(10) => next_NPC_10_port, 
                           DATA_IN(9) => next_NPC_9_port, DATA_IN(8) => 
                           next_NPC_8_port, DATA_IN(7) => next_NPC_7_port, 
                           DATA_IN(6) => next_NPC_6_port, DATA_IN(5) => 
                           next_NPC_5_port, DATA_IN(4) => next_NPC_4_port, 
                           DATA_IN(3) => next_NPC_3_port, DATA_IN(2) => 
                           next_NPC_2_port, DATA_IN(1) => next_NPC_1_port, 
                           DATA_IN(0) => next_NPC_0_port, DATA_OUT(31) => 
                           current_NPC_31_port, DATA_OUT(30) => 
                           current_NPC_30_port, DATA_OUT(29) => 
                           current_NPC_29_port, DATA_OUT(28) => 
                           current_NPC_28_port, DATA_OUT(27) => 
                           current_NPC_27_port, DATA_OUT(26) => 
                           current_NPC_26_port, DATA_OUT(25) => 
                           current_NPC_25_port, DATA_OUT(24) => 
                           current_NPC_24_port, DATA_OUT(23) => 
                           current_NPC_23_port, DATA_OUT(22) => 
                           current_NPC_22_port, DATA_OUT(21) => 
                           current_NPC_21_port, DATA_OUT(20) => 
                           current_NPC_20_port, DATA_OUT(19) => 
                           current_NPC_19_port, DATA_OUT(18) => 
                           current_NPC_18_port, DATA_OUT(17) => 
                           current_NPC_17_port, DATA_OUT(16) => 
                           current_NPC_16_port, DATA_OUT(15) => 
                           current_NPC_15_port, DATA_OUT(14) => 
                           current_NPC_14_port, DATA_OUT(13) => 
                           current_NPC_13_port, DATA_OUT(12) => 
                           current_NPC_12_port, DATA_OUT(11) => 
                           current_NPC_11_port, DATA_OUT(10) => 
                           current_NPC_10_port, DATA_OUT(9) => 
                           current_NPC_9_port, DATA_OUT(8) => 
                           current_NPC_8_port, DATA_OUT(7) => 
                           current_NPC_7_port, DATA_OUT(6) => 
                           current_NPC_6_port, DATA_OUT(5) => 
                           current_NPC_5_port, DATA_OUT(4) => 
                           current_NPC_4_port, DATA_OUT(3) => 
                           current_NPC_3_port, DATA_OUT(2) => 
                           current_NPC_2_port, DATA_OUT(1) => 
                           current_NPC_1_port, DATA_OUT(0) => 
                           current_NPC_0_port);
   IR_REG : REG_GENERIC_NBIT32_4 port map( CLK => CLK, RST => RST, EN => 
                           IR_LATCH_EN, DATA_IN(31) => IR_IN(31), DATA_IN(30) 
                           => IR_IN(30), DATA_IN(29) => IR_IN(29), DATA_IN(28) 
                           => IR_IN(28), DATA_IN(27) => IR_IN(27), DATA_IN(26) 
                           => IR_IN(26), DATA_IN(25) => IR_IN(25), DATA_IN(24) 
                           => IR_IN(24), DATA_IN(23) => IR_IN(23), DATA_IN(22) 
                           => IR_IN(22), DATA_IN(21) => IR_IN(21), DATA_IN(20) 
                           => IR_IN(20), DATA_IN(19) => IR_IN(19), DATA_IN(18) 
                           => IR_IN(18), DATA_IN(17) => IR_IN(17), DATA_IN(16) 
                           => IR_IN(16), DATA_IN(15) => IR_IN(15), DATA_IN(14) 
                           => IR_IN(14), DATA_IN(13) => IR_IN(13), DATA_IN(12) 
                           => IR_IN(12), DATA_IN(11) => IR_IN(11), DATA_IN(10) 
                           => IR_IN(10), DATA_IN(9) => IR_IN(9), DATA_IN(8) => 
                           IR_IN(8), DATA_IN(7) => IR_IN(7), DATA_IN(6) => 
                           IR_IN(6), DATA_IN(5) => IR_IN(5), DATA_IN(4) => 
                           IR_IN(4), DATA_IN(3) => IR_IN(3), DATA_IN(2) => 
                           IR_IN(2), DATA_IN(1) => IR_IN(1), DATA_IN(0) => 
                           IR_IN(0), DATA_OUT(31) => n_1607, DATA_OUT(30) => 
                           n_1608, DATA_OUT(29) => n_1609, DATA_OUT(28) => 
                           n_1610, DATA_OUT(27) => n_1611, DATA_OUT(26) => 
                           n_1612, DATA_OUT(25) => current_IW_25_port, 
                           DATA_OUT(24) => current_IW_24_port, DATA_OUT(23) => 
                           current_IW_23_port, DATA_OUT(22) => 
                           current_IW_22_port, DATA_OUT(21) => 
                           current_IW_21_port, DATA_OUT(20) => 
                           current_IW_20_port, DATA_OUT(19) => 
                           current_IW_19_port, DATA_OUT(18) => 
                           current_IW_18_port, DATA_OUT(17) => 
                           current_IW_17_port, DATA_OUT(16) => 
                           current_IW_16_port, DATA_OUT(15) => 
                           current_IW_15_port, DATA_OUT(14) => 
                           current_IW_14_port, DATA_OUT(13) => 
                           current_IW_13_port, DATA_OUT(12) => 
                           current_IW_12_port, DATA_OUT(11) => 
                           current_IW_11_port, DATA_OUT(10) => 
                           current_IW_10_port, DATA_OUT(9) => current_IW_9_port
                           , DATA_OUT(8) => current_IW_8_port, DATA_OUT(7) => 
                           current_IW_7_port, DATA_OUT(6) => current_IW_6_port,
                           DATA_OUT(5) => current_IW_5_port, DATA_OUT(4) => 
                           current_IW_4_port, DATA_OUT(3) => current_IW_3_port,
                           DATA_OUT(2) => current_IW_2_port, DATA_OUT(1) => 
                           current_IW_1_port, DATA_OUT(0) => current_IW_0_port)
                           ;
   IMM_REG : REG_GENERIC_NBIT26 port map( CLK => CLK, RST => RST, EN => 
                           RegIMM_LATCH_EN, DATA_IN(25) => current_IW_25_port, 
                           DATA_IN(24) => current_IW_24_port, DATA_IN(23) => 
                           current_IW_23_port, DATA_IN(22) => 
                           current_IW_22_port, DATA_IN(21) => 
                           current_IW_21_port, DATA_IN(20) => 
                           current_IW_20_port, DATA_IN(19) => 
                           current_IW_19_port, DATA_IN(18) => 
                           current_IW_18_port, DATA_IN(17) => 
                           current_IW_17_port, DATA_IN(16) => 
                           current_IW_16_port, DATA_IN(15) => 
                           current_IW_15_port, DATA_IN(14) => 
                           current_IW_14_port, DATA_IN(13) => 
                           current_IW_13_port, DATA_IN(12) => 
                           current_IW_12_port, DATA_IN(11) => 
                           current_IW_11_port, DATA_IN(10) => 
                           current_IW_10_port, DATA_IN(9) => current_IW_9_port,
                           DATA_IN(8) => current_IW_8_port, DATA_IN(7) => 
                           current_IW_7_port, DATA_IN(6) => current_IW_6_port, 
                           DATA_IN(5) => current_IW_5_port, DATA_IN(4) => 
                           current_IW_4_port, DATA_IN(3) => current_IW_3_port, 
                           DATA_IN(2) => current_IW_2_port, DATA_IN(1) => 
                           current_IW_1_port, DATA_IN(0) => current_IW_0_port, 
                           DATA_OUT(25) => IMM_IN_25_port, DATA_OUT(24) => 
                           IMM_IN_24_port, DATA_OUT(23) => IMM_IN_23_port, 
                           DATA_OUT(22) => IMM_IN_22_port, DATA_OUT(21) => 
                           IMM_IN_21_port, DATA_OUT(20) => IMM_IN_20_port, 
                           DATA_OUT(19) => IMM_IN_19_port, DATA_OUT(18) => 
                           IMM_IN_18_port, DATA_OUT(17) => IMM_IN_17_port, 
                           DATA_OUT(16) => IMM_IN_16_port, DATA_OUT(15) => 
                           IMM_IN_15_port, DATA_OUT(14) => IMM_IN_14_port, 
                           DATA_OUT(13) => IMM_IN_13_port, DATA_OUT(12) => 
                           IMM_IN_12_port, DATA_OUT(11) => IMM_IN_11_port, 
                           DATA_OUT(10) => IMM_IN_10_port, DATA_OUT(9) => 
                           IMM_IN_9_port, DATA_OUT(8) => IMM_IN_8_port, 
                           DATA_OUT(7) => IMM_IN_7_port, DATA_OUT(6) => 
                           IMM_IN_6_port, DATA_OUT(5) => IMM_IN_5_port, 
                           DATA_OUT(4) => IMM_IN_4_port, DATA_OUT(3) => 
                           IMM_IN_3_port, DATA_OUT(2) => IMM_IN_2_port, 
                           DATA_OUT(1) => IMM_IN_1_port, DATA_OUT(0) => 
                           IMM_IN_0_port);
   WB1_REG : REG_GENERIC_NBIT5_0 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, DATA_IN(4) => WB1_IN_4_port, 
                           DATA_IN(3) => WB1_IN_3_port, DATA_IN(2) => 
                           WB1_IN_2_port, DATA_IN(1) => WB1_IN_1_port, 
                           DATA_IN(0) => WB1_IN_0_port, DATA_OUT(4) => 
                           WB2_IN_4_port, DATA_OUT(3) => WB2_IN_3_port, 
                           DATA_OUT(2) => WB2_IN_2_port, DATA_OUT(1) => 
                           WB2_IN_1_port, DATA_OUT(0) => WB2_IN_0_port);
   WB2_REG : REG_GENERIC_NBIT5_2 port map( CLK => CLK, RST => RST, EN => 
                           ALU_OUTREG_EN, DATA_IN(4) => WB2_IN_4_port, 
                           DATA_IN(3) => WB2_IN_3_port, DATA_IN(2) => 
                           WB2_IN_2_port, DATA_IN(1) => WB2_IN_1_port, 
                           DATA_IN(0) => WB2_IN_0_port, DATA_OUT(4) => 
                           WB2_OUT_4_port, DATA_OUT(3) => WB2_OUT_3_port, 
                           DATA_OUT(2) => WB2_OUT_2_port, DATA_OUT(1) => 
                           WB2_OUT_1_port, DATA_OUT(0) => WB2_OUT_0_port);
   WB3_REG : REG_GENERIC_NBIT5_1 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, DATA_IN(4) => WB2_OUT_4_port, 
                           DATA_IN(3) => WB2_OUT_3_port, DATA_IN(2) => 
                           WB2_OUT_2_port, DATA_IN(1) => WB2_OUT_1_port, 
                           DATA_IN(0) => WB2_OUT_0_port, DATA_OUT(4) => 
                           WB3_OUT_4_port, DATA_OUT(3) => WB3_OUT_3_port, 
                           DATA_OUT(2) => WB3_OUT_2_port, DATA_OUT(1) => 
                           WB3_OUT_1_port, DATA_OUT(0) => WB3_OUT_0_port);
   ALU_OUT_REG : REG_GENERIC_NBIT32_3 port map( CLK => CLK, RST => RST, EN => 
                           ALU_OUTREG_EN, DATA_IN(31) => next_ALU_OUT_31_port, 
                           DATA_IN(30) => next_ALU_OUT_30_port, DATA_IN(29) => 
                           next_ALU_OUT_29_port, DATA_IN(28) => 
                           next_ALU_OUT_28_port, DATA_IN(27) => 
                           next_ALU_OUT_27_port, DATA_IN(26) => 
                           next_ALU_OUT_26_port, DATA_IN(25) => 
                           next_ALU_OUT_25_port, DATA_IN(24) => 
                           next_ALU_OUT_24_port, DATA_IN(23) => 
                           next_ALU_OUT_23_port, DATA_IN(22) => 
                           next_ALU_OUT_22_port, DATA_IN(21) => 
                           next_ALU_OUT_21_port, DATA_IN(20) => 
                           next_ALU_OUT_20_port, DATA_IN(19) => 
                           next_ALU_OUT_19_port, DATA_IN(18) => 
                           next_ALU_OUT_18_port, DATA_IN(17) => 
                           next_ALU_OUT_17_port, DATA_IN(16) => 
                           next_ALU_OUT_16_port, DATA_IN(15) => 
                           next_ALU_OUT_15_port, DATA_IN(14) => 
                           next_ALU_OUT_14_port, DATA_IN(13) => 
                           next_ALU_OUT_13_port, DATA_IN(12) => 
                           next_ALU_OUT_12_port, DATA_IN(11) => 
                           next_ALU_OUT_11_port, DATA_IN(10) => 
                           next_ALU_OUT_10_port, DATA_IN(9) => 
                           next_ALU_OUT_9_port, DATA_IN(8) => 
                           next_ALU_OUT_8_port, DATA_IN(7) => 
                           next_ALU_OUT_7_port, DATA_IN(6) => 
                           next_ALU_OUT_6_port, DATA_IN(5) => 
                           next_ALU_OUT_5_port, DATA_IN(4) => 
                           next_ALU_OUT_4_port, DATA_IN(3) => 
                           next_ALU_OUT_3_port, DATA_IN(2) => 
                           next_ALU_OUT_2_port, DATA_IN(1) => 
                           next_ALU_OUT_1_port, DATA_IN(0) => 
                           next_ALU_OUT_0_port, DATA_OUT(31) => 
                           current_ALU_OUT_31_port, DATA_OUT(30) => 
                           current_ALU_OUT_30_port, DATA_OUT(29) => 
                           current_ALU_OUT_29_port, DATA_OUT(28) => 
                           current_ALU_OUT_28_port, DATA_OUT(27) => 
                           current_ALU_OUT_27_port, DATA_OUT(26) => 
                           current_ALU_OUT_26_port, DATA_OUT(25) => 
                           current_ALU_OUT_25_port, DATA_OUT(24) => 
                           current_ALU_OUT_24_port, DATA_OUT(23) => 
                           current_ALU_OUT_23_port, DATA_OUT(22) => 
                           current_ALU_OUT_22_port, DATA_OUT(21) => 
                           current_ALU_OUT_21_port, DATA_OUT(20) => 
                           current_ALU_OUT_20_port, DATA_OUT(19) => 
                           current_ALU_OUT_19_port, DATA_OUT(18) => 
                           current_ALU_OUT_18_port, DATA_OUT(17) => 
                           current_ALU_OUT_17_port, DATA_OUT(16) => 
                           current_ALU_OUT_16_port, DATA_OUT(15) => 
                           current_ALU_OUT_15_port, DATA_OUT(14) => 
                           current_ALU_OUT_14_port, DATA_OUT(13) => 
                           current_ALU_OUT_13_port, DATA_OUT(12) => 
                           current_ALU_OUT_12_port, DATA_OUT(11) => 
                           current_ALU_OUT_11_port, DATA_OUT(10) => 
                           current_ALU_OUT_10_port, DATA_OUT(9) => 
                           current_ALU_OUT_9_port, DATA_OUT(8) => 
                           current_ALU_OUT_8_port, DATA_OUT(7) => 
                           current_ALU_OUT_7_port, DATA_OUT(6) => 
                           current_ALU_OUT_6_port, DATA_OUT(5) => D_ADDR_5_port
                           , DATA_OUT(4) => D_ADDR_4_port, DATA_OUT(3) => 
                           D_ADDR_3_port, DATA_OUT(2) => D_ADDR_2_port, 
                           DATA_OUT(1) => D_ADDR_1_port, DATA_OUT(0) => 
                           D_ADDR_0_port);
   B_OUT_REG : REG_GENERIC_NBIT32_2 port map( CLK => CLK, RST => RST, EN => 
                           ALU_OUTREG_EN, DATA_IN(31) => B_OUT_31_port, 
                           DATA_IN(30) => B_OUT_30_port, DATA_IN(29) => 
                           B_OUT_29_port, DATA_IN(28) => B_OUT_28_port, 
                           DATA_IN(27) => B_OUT_27_port, DATA_IN(26) => 
                           B_OUT_26_port, DATA_IN(25) => B_OUT_25_port, 
                           DATA_IN(24) => B_OUT_24_port, DATA_IN(23) => 
                           B_OUT_23_port, DATA_IN(22) => B_OUT_22_port, 
                           DATA_IN(21) => B_OUT_21_port, DATA_IN(20) => 
                           B_OUT_20_port, DATA_IN(19) => B_OUT_19_port, 
                           DATA_IN(18) => B_OUT_18_port, DATA_IN(17) => 
                           B_OUT_17_port, DATA_IN(16) => B_OUT_16_port, 
                           DATA_IN(15) => B_OUT_15_port, DATA_IN(14) => 
                           B_OUT_14_port, DATA_IN(13) => B_OUT_13_port, 
                           DATA_IN(12) => B_OUT_12_port, DATA_IN(11) => 
                           B_OUT_11_port, DATA_IN(10) => B_OUT_10_port, 
                           DATA_IN(9) => B_OUT_9_port, DATA_IN(8) => 
                           B_OUT_8_port, DATA_IN(7) => B_OUT_7_port, DATA_IN(6)
                           => B_OUT_6_port, DATA_IN(5) => B_OUT_5_port, 
                           DATA_IN(4) => B_OUT_4_port, DATA_IN(3) => 
                           B_OUT_3_port, DATA_IN(2) => B_OUT_2_port, DATA_IN(1)
                           => B_OUT_1_port, DATA_IN(0) => B_OUT_0_port, 
                           DATA_OUT(31) => D_DATA_IN(31), DATA_OUT(30) => 
                           D_DATA_IN(30), DATA_OUT(29) => D_DATA_IN(29), 
                           DATA_OUT(28) => D_DATA_IN(28), DATA_OUT(27) => 
                           D_DATA_IN(27), DATA_OUT(26) => D_DATA_IN(26), 
                           DATA_OUT(25) => D_DATA_IN(25), DATA_OUT(24) => 
                           D_DATA_IN(24), DATA_OUT(23) => D_DATA_IN(23), 
                           DATA_OUT(22) => D_DATA_IN(22), DATA_OUT(21) => 
                           D_DATA_IN(21), DATA_OUT(20) => D_DATA_IN(20), 
                           DATA_OUT(19) => D_DATA_IN(19), DATA_OUT(18) => 
                           D_DATA_IN(18), DATA_OUT(17) => D_DATA_IN(17), 
                           DATA_OUT(16) => D_DATA_IN(16), DATA_OUT(15) => 
                           D_DATA_IN(15), DATA_OUT(14) => D_DATA_IN(14), 
                           DATA_OUT(13) => D_DATA_IN(13), DATA_OUT(12) => 
                           D_DATA_IN(12), DATA_OUT(11) => D_DATA_IN(11), 
                           DATA_OUT(10) => D_DATA_IN(10), DATA_OUT(9) => 
                           D_DATA_IN(9), DATA_OUT(8) => D_DATA_IN(8), 
                           DATA_OUT(7) => D_DATA_IN(7), DATA_OUT(6) => 
                           D_DATA_IN(6), DATA_OUT(5) => D_DATA_IN(5), 
                           DATA_OUT(4) => D_DATA_IN(4), DATA_OUT(3) => 
                           D_DATA_IN(3), DATA_OUT(2) => D_DATA_IN(2), 
                           DATA_OUT(1) => D_DATA_IN(1), DATA_OUT(0) => 
                           D_DATA_IN(0));
   ALU_OUT_REG2 : REG_GENERIC_NBIT32_1 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, DATA_IN(31) => 
                           current_ALU_OUT_31_port, DATA_IN(30) => 
                           current_ALU_OUT_30_port, DATA_IN(29) => 
                           current_ALU_OUT_29_port, DATA_IN(28) => 
                           current_ALU_OUT_28_port, DATA_IN(27) => 
                           current_ALU_OUT_27_port, DATA_IN(26) => 
                           current_ALU_OUT_26_port, DATA_IN(25) => 
                           current_ALU_OUT_25_port, DATA_IN(24) => 
                           current_ALU_OUT_24_port, DATA_IN(23) => 
                           current_ALU_OUT_23_port, DATA_IN(22) => 
                           current_ALU_OUT_22_port, DATA_IN(21) => 
                           current_ALU_OUT_21_port, DATA_IN(20) => 
                           current_ALU_OUT_20_port, DATA_IN(19) => 
                           current_ALU_OUT_19_port, DATA_IN(18) => 
                           current_ALU_OUT_18_port, DATA_IN(17) => 
                           current_ALU_OUT_17_port, DATA_IN(16) => 
                           current_ALU_OUT_16_port, DATA_IN(15) => 
                           current_ALU_OUT_15_port, DATA_IN(14) => 
                           current_ALU_OUT_14_port, DATA_IN(13) => 
                           current_ALU_OUT_13_port, DATA_IN(12) => 
                           current_ALU_OUT_12_port, DATA_IN(11) => 
                           current_ALU_OUT_11_port, DATA_IN(10) => 
                           current_ALU_OUT_10_port, DATA_IN(9) => 
                           current_ALU_OUT_9_port, DATA_IN(8) => 
                           current_ALU_OUT_8_port, DATA_IN(7) => 
                           current_ALU_OUT_7_port, DATA_IN(6) => 
                           current_ALU_OUT_6_port, DATA_IN(5) => D_ADDR_5_port,
                           DATA_IN(4) => D_ADDR_4_port, DATA_IN(3) => 
                           D_ADDR_3_port, DATA_IN(2) => D_ADDR_2_port, 
                           DATA_IN(1) => D_ADDR_1_port, DATA_IN(0) => 
                           D_ADDR_0_port, DATA_OUT(31) => 
                           current_ALU_OUT2_31_port, DATA_OUT(30) => 
                           current_ALU_OUT2_30_port, DATA_OUT(29) => 
                           current_ALU_OUT2_29_port, DATA_OUT(28) => 
                           current_ALU_OUT2_28_port, DATA_OUT(27) => 
                           current_ALU_OUT2_27_port, DATA_OUT(26) => 
                           current_ALU_OUT2_26_port, DATA_OUT(25) => 
                           current_ALU_OUT2_25_port, DATA_OUT(24) => 
                           current_ALU_OUT2_24_port, DATA_OUT(23) => 
                           current_ALU_OUT2_23_port, DATA_OUT(22) => 
                           current_ALU_OUT2_22_port, DATA_OUT(21) => 
                           current_ALU_OUT2_21_port, DATA_OUT(20) => 
                           current_ALU_OUT2_20_port, DATA_OUT(19) => 
                           current_ALU_OUT2_19_port, DATA_OUT(18) => 
                           current_ALU_OUT2_18_port, DATA_OUT(17) => 
                           current_ALU_OUT2_17_port, DATA_OUT(16) => 
                           current_ALU_OUT2_16_port, DATA_OUT(15) => 
                           current_ALU_OUT2_15_port, DATA_OUT(14) => 
                           current_ALU_OUT2_14_port, DATA_OUT(13) => 
                           current_ALU_OUT2_13_port, DATA_OUT(12) => 
                           current_ALU_OUT2_12_port, DATA_OUT(11) => 
                           current_ALU_OUT2_11_port, DATA_OUT(10) => 
                           current_ALU_OUT2_10_port, DATA_OUT(9) => 
                           current_ALU_OUT2_9_port, DATA_OUT(8) => 
                           current_ALU_OUT2_8_port, DATA_OUT(7) => 
                           current_ALU_OUT2_7_port, DATA_OUT(6) => 
                           current_ALU_OUT2_6_port, DATA_OUT(5) => 
                           current_ALU_OUT2_5_port, DATA_OUT(4) => 
                           current_ALU_OUT2_4_port, DATA_OUT(3) => 
                           current_ALU_OUT2_3_port, DATA_OUT(2) => 
                           current_ALU_OUT2_2_port, DATA_OUT(1) => 
                           current_ALU_OUT2_1_port, DATA_OUT(0) => 
                           current_ALU_OUT2_0_port);
   BU : BRANCHING_UNIT_N32 port map( CLK => CLK, RST => RST, Reg_A(31) => 
                           A_OUT_31_port, Reg_A(30) => A_OUT_30_port, Reg_A(29)
                           => A_OUT_29_port, Reg_A(28) => A_OUT_28_port, 
                           Reg_A(27) => A_OUT_27_port, Reg_A(26) => 
                           A_OUT_26_port, Reg_A(25) => A_OUT_25_port, Reg_A(24)
                           => A_OUT_24_port, Reg_A(23) => A_OUT_23_port, 
                           Reg_A(22) => A_OUT_22_port, Reg_A(21) => 
                           A_OUT_21_port, Reg_A(20) => A_OUT_20_port, Reg_A(19)
                           => A_OUT_19_port, Reg_A(18) => A_OUT_18_port, 
                           Reg_A(17) => A_OUT_17_port, Reg_A(16) => 
                           A_OUT_16_port, Reg_A(15) => A_OUT_15_port, Reg_A(14)
                           => A_OUT_14_port, Reg_A(13) => A_OUT_13_port, 
                           Reg_A(12) => A_OUT_12_port, Reg_A(11) => 
                           A_OUT_11_port, Reg_A(10) => A_OUT_10_port, Reg_A(9) 
                           => A_OUT_9_port, Reg_A(8) => A_OUT_8_port, Reg_A(7) 
                           => A_OUT_7_port, Reg_A(6) => A_OUT_6_port, Reg_A(5) 
                           => A_OUT_5_port, Reg_A(4) => A_OUT_4_port, Reg_A(3) 
                           => A_OUT_3_port, Reg_A(2) => A_OUT_2_port, Reg_A(1) 
                           => A_OUT_1_port, Reg_A(0) => A_OUT_0_port, EQ_cond 
                           => EQ_COND, IS_JUMP => IS_JUMP, branch_taken => 
                           branch_taken);
   PC_MUX : MUX21_GENERIC_NBIT32_0 port map( A(31) => current_NPC_31_port, 
                           A(30) => current_NPC_30_port, A(29) => 
                           current_NPC_29_port, A(28) => current_NPC_28_port, 
                           A(27) => current_NPC_27_port, A(26) => 
                           current_NPC_26_port, A(25) => current_NPC_25_port, 
                           A(24) => current_NPC_24_port, A(23) => 
                           current_NPC_23_port, A(22) => current_NPC_22_port, 
                           A(21) => current_NPC_21_port, A(20) => 
                           current_NPC_20_port, A(19) => current_NPC_19_port, 
                           A(18) => current_NPC_18_port, A(17) => 
                           current_NPC_17_port, A(16) => current_NPC_16_port, 
                           A(15) => current_NPC_15_port, A(14) => 
                           current_NPC_14_port, A(13) => current_NPC_13_port, 
                           A(12) => current_NPC_12_port, A(11) => 
                           current_NPC_11_port, A(10) => current_NPC_10_port, 
                           A(9) => current_NPC_9_port, A(8) => 
                           current_NPC_8_port, A(7) => current_NPC_7_port, A(6)
                           => current_NPC_6_port, A(5) => current_NPC_5_port, 
                           A(4) => current_NPC_4_port, A(3) => 
                           current_NPC_3_port, A(2) => current_NPC_2_port, A(1)
                           => current_NPC_1_port, A(0) => current_NPC_0_port, 
                           B(31) => current_ALU_OUT_31_port, B(30) => 
                           current_ALU_OUT_30_port, B(29) => 
                           current_ALU_OUT_29_port, B(28) => 
                           current_ALU_OUT_28_port, B(27) => 
                           current_ALU_OUT_27_port, B(26) => 
                           current_ALU_OUT_26_port, B(25) => 
                           current_ALU_OUT_25_port, B(24) => 
                           current_ALU_OUT_24_port, B(23) => 
                           current_ALU_OUT_23_port, B(22) => 
                           current_ALU_OUT_22_port, B(21) => 
                           current_ALU_OUT_21_port, B(20) => 
                           current_ALU_OUT_20_port, B(19) => 
                           current_ALU_OUT_19_port, B(18) => 
                           current_ALU_OUT_18_port, B(17) => 
                           current_ALU_OUT_17_port, B(16) => 
                           current_ALU_OUT_16_port, B(15) => 
                           current_ALU_OUT_15_port, B(14) => 
                           current_ALU_OUT_14_port, B(13) => 
                           current_ALU_OUT_13_port, B(12) => 
                           current_ALU_OUT_12_port, B(11) => 
                           current_ALU_OUT_11_port, B(10) => 
                           current_ALU_OUT_10_port, B(9) => 
                           current_ALU_OUT_9_port, B(8) => 
                           current_ALU_OUT_8_port, B(7) => 
                           current_ALU_OUT_7_port, B(6) => 
                           current_ALU_OUT_6_port, B(5) => D_ADDR_5_port, B(4) 
                           => D_ADDR_4_port, B(3) => D_ADDR_3_port, B(2) => 
                           D_ADDR_2_port, B(1) => D_ADDR_1_port, B(0) => 
                           D_ADDR_0_port, SEL => PC_MUX_SEL, Y(31) => 
                           PC_BUS_31_port, Y(30) => PC_BUS_30_port, Y(29) => 
                           PC_BUS_29_port, Y(28) => PC_BUS_28_port, Y(27) => 
                           PC_BUS_27_port, Y(26) => PC_BUS_26_port, Y(25) => 
                           PC_BUS_25_port, Y(24) => PC_BUS_24_port, Y(23) => 
                           PC_BUS_23_port, Y(22) => PC_BUS_22_port, Y(21) => 
                           PC_BUS_21_port, Y(20) => PC_BUS_20_port, Y(19) => 
                           PC_BUS_19_port, Y(18) => PC_BUS_18_port, Y(17) => 
                           PC_BUS_17_port, Y(16) => PC_BUS_16_port, Y(15) => 
                           PC_BUS_15_port, Y(14) => PC_BUS_14_port, Y(13) => 
                           PC_BUS_13_port, Y(12) => PC_BUS_12_port, Y(11) => 
                           PC_BUS_11_port, Y(10) => PC_BUS_10_port, Y(9) => 
                           PC_BUS_9_port, Y(8) => PC_BUS_8_port, Y(7) => 
                           PC_BUS_7_port, Y(6) => PC_BUS_6_port, Y(5) => 
                           PC_BUS_5_port, Y(4) => PC_BUS_4_port, Y(3) => 
                           PC_BUS_3_port, Y(2) => PC_BUS_2_port, Y(1) => 
                           PC_BUS_1_port, Y(0) => PC_BUS_0_port);
   J_MUX : MUX21 port map( A => X_Logic0_port, B => branch_taken, SEL => 
                           JUMP_EN, Y => PC_MUX_SEL);
   RD_MUX : MUX21_GENERIC_NBIT5_0 port map( A(4) => current_IW_15_port, A(3) =>
                           current_IW_14_port, A(2) => current_IW_13_port, A(1)
                           => current_IW_12_port, A(0) => current_IW_11_port, 
                           B(4) => current_IW_20_port, B(3) => 
                           current_IW_19_port, B(2) => current_IW_18_port, B(1)
                           => current_IW_17_port, B(0) => current_IW_16_port, 
                           SEL => RegIMM_LATCH_EN, Y(4) => WB1_IN_4_port, Y(3) 
                           => WB1_IN_3_port, Y(2) => WB1_IN_2_port, Y(1) => 
                           WB1_IN_1_port, Y(0) => WB1_IN_0_port);
   OP1_MUX : MUX21_GENERIC_NBIT32_4 port map( A(31) => A_OUT_31_port, A(30) => 
                           A_OUT_30_port, A(29) => A_OUT_29_port, A(28) => 
                           A_OUT_28_port, A(27) => A_OUT_27_port, A(26) => 
                           A_OUT_26_port, A(25) => A_OUT_25_port, A(24) => 
                           A_OUT_24_port, A(23) => A_OUT_23_port, A(22) => 
                           A_OUT_22_port, A(21) => A_OUT_21_port, A(20) => 
                           A_OUT_20_port, A(19) => A_OUT_19_port, A(18) => 
                           A_OUT_18_port, A(17) => A_OUT_17_port, A(16) => 
                           A_OUT_16_port, A(15) => A_OUT_15_port, A(14) => 
                           A_OUT_14_port, A(13) => A_OUT_13_port, A(12) => 
                           A_OUT_12_port, A(11) => A_OUT_11_port, A(10) => 
                           A_OUT_10_port, A(9) => A_OUT_9_port, A(8) => 
                           A_OUT_8_port, A(7) => A_OUT_7_port, A(6) => 
                           A_OUT_6_port, A(5) => A_OUT_5_port, A(4) => 
                           A_OUT_4_port, A(3) => A_OUT_3_port, A(2) => 
                           A_OUT_2_port, A(1) => A_OUT_1_port, A(0) => 
                           A_OUT_0_port, B(31) => current_PC1_31_port, B(30) =>
                           current_PC1_30_port, B(29) => current_PC1_29_port, 
                           B(28) => current_PC1_28_port, B(27) => 
                           current_PC1_27_port, B(26) => current_PC1_26_port, 
                           B(25) => current_PC1_25_port, B(24) => 
                           current_PC1_24_port, B(23) => current_PC1_23_port, 
                           B(22) => current_PC1_22_port, B(21) => 
                           current_PC1_21_port, B(20) => current_PC1_20_port, 
                           B(19) => current_PC1_19_port, B(18) => 
                           current_PC1_18_port, B(17) => current_PC1_17_port, 
                           B(16) => current_PC1_16_port, B(15) => 
                           current_PC1_15_port, B(14) => current_PC1_14_port, 
                           B(13) => current_PC1_13_port, B(12) => 
                           current_PC1_12_port, B(11) => current_PC1_11_port, 
                           B(10) => current_PC1_10_port, B(9) => 
                           current_PC1_9_port, B(8) => current_PC1_8_port, B(7)
                           => current_PC1_7_port, B(6) => current_PC1_6_port, 
                           B(5) => current_PC1_5_port, B(4) => 
                           current_PC1_4_port, B(3) => current_PC1_3_port, B(2)
                           => current_PC1_2_port, B(1) => current_PC1_1_port, 
                           B(0) => current_PC1_0_port, SEL => MUXA_SEL, Y(31) 
                           => ALU_OP1_31_port, Y(30) => ALU_OP1_30_port, Y(29) 
                           => ALU_OP1_29_port, Y(28) => ALU_OP1_28_port, Y(27) 
                           => ALU_OP1_27_port, Y(26) => ALU_OP1_26_port, Y(25) 
                           => ALU_OP1_25_port, Y(24) => ALU_OP1_24_port, Y(23) 
                           => ALU_OP1_23_port, Y(22) => ALU_OP1_22_port, Y(21) 
                           => ALU_OP1_21_port, Y(20) => ALU_OP1_20_port, Y(19) 
                           => ALU_OP1_19_port, Y(18) => ALU_OP1_18_port, Y(17) 
                           => ALU_OP1_17_port, Y(16) => ALU_OP1_16_port, Y(15) 
                           => ALU_OP1_15_port, Y(14) => ALU_OP1_14_port, Y(13) 
                           => ALU_OP1_13_port, Y(12) => ALU_OP1_12_port, Y(11) 
                           => ALU_OP1_11_port, Y(10) => ALU_OP1_10_port, Y(9) 
                           => ALU_OP1_9_port, Y(8) => ALU_OP1_8_port, Y(7) => 
                           ALU_OP1_7_port, Y(6) => ALU_OP1_6_port, Y(5) => 
                           ALU_OP1_5_port, Y(4) => ALU_OP1_4_port, Y(3) => 
                           ALU_OP1_3_port, Y(2) => ALU_OP1_2_port, Y(1) => 
                           ALU_OP1_1_port, Y(0) => ALU_OP1_0_port);
   OP2_MUX : MUX21_GENERIC_NBIT32_3 port map( A(31) => B_OUT_31_port, A(30) => 
                           B_OUT_30_port, A(29) => B_OUT_29_port, A(28) => 
                           B_OUT_28_port, A(27) => B_OUT_27_port, A(26) => 
                           B_OUT_26_port, A(25) => B_OUT_25_port, A(24) => 
                           B_OUT_24_port, A(23) => B_OUT_23_port, A(22) => 
                           B_OUT_22_port, A(21) => B_OUT_21_port, A(20) => 
                           B_OUT_20_port, A(19) => B_OUT_19_port, A(18) => 
                           B_OUT_18_port, A(17) => B_OUT_17_port, A(16) => 
                           B_OUT_16_port, A(15) => B_OUT_15_port, A(14) => 
                           B_OUT_14_port, A(13) => B_OUT_13_port, A(12) => 
                           B_OUT_12_port, A(11) => B_OUT_11_port, A(10) => 
                           B_OUT_10_port, A(9) => B_OUT_9_port, A(8) => 
                           B_OUT_8_port, A(7) => B_OUT_7_port, A(6) => 
                           B_OUT_6_port, A(5) => B_OUT_5_port, A(4) => 
                           B_OUT_4_port, A(3) => B_OUT_3_port, A(2) => 
                           B_OUT_2_port, A(1) => B_OUT_1_port, A(0) => 
                           B_OUT_0_port, B(31) => IMM_OUT_31_port, B(30) => 
                           IMM_OUT_30_port, B(29) => IMM_OUT_29_port, B(28) => 
                           IMM_OUT_28_port, B(27) => IMM_OUT_27_port, B(26) => 
                           IMM_OUT_26_port, B(25) => IMM_OUT_25_port, B(24) => 
                           IMM_OUT_24_port, B(23) => IMM_OUT_23_port, B(22) => 
                           IMM_OUT_22_port, B(21) => IMM_OUT_21_port, B(20) => 
                           IMM_OUT_20_port, B(19) => IMM_OUT_19_port, B(18) => 
                           IMM_OUT_18_port, B(17) => IMM_OUT_17_port, B(16) => 
                           IMM_OUT_16_port, B(15) => IMM_OUT_15_port, B(14) => 
                           IMM_OUT_14_port, B(13) => IMM_OUT_13_port, B(12) => 
                           IMM_OUT_12_port, B(11) => IMM_OUT_11_port, B(10) => 
                           IMM_OUT_10_port, B(9) => IMM_OUT_9_port, B(8) => 
                           IMM_OUT_8_port, B(7) => IMM_OUT_7_port, B(6) => 
                           IMM_OUT_6_port, B(5) => IMM_OUT_5_port, B(4) => 
                           IMM_OUT_4_port, B(3) => IMM_OUT_3_port, B(2) => 
                           IMM_OUT_2_port, B(1) => IMM_OUT_1_port, B(0) => 
                           IMM_OUT_0_port, SEL => MUXB_SEL, Y(31) => 
                           ALU_OP2_31_port, Y(30) => ALU_OP2_30_port, Y(29) => 
                           ALU_OP2_29_port, Y(28) => ALU_OP2_28_port, Y(27) => 
                           ALU_OP2_27_port, Y(26) => ALU_OP2_26_port, Y(25) => 
                           ALU_OP2_25_port, Y(24) => ALU_OP2_24_port, Y(23) => 
                           ALU_OP2_23_port, Y(22) => ALU_OP2_22_port, Y(21) => 
                           ALU_OP2_21_port, Y(20) => ALU_OP2_20_port, Y(19) => 
                           ALU_OP2_19_port, Y(18) => ALU_OP2_18_port, Y(17) => 
                           ALU_OP2_17_port, Y(16) => ALU_OP2_16_port, Y(15) => 
                           ALU_OP2_15_port, Y(14) => ALU_OP2_14_port, Y(13) => 
                           ALU_OP2_13_port, Y(12) => ALU_OP2_12_port, Y(11) => 
                           ALU_OP2_11_port, Y(10) => ALU_OP2_10_port, Y(9) => 
                           ALU_OP2_9_port, Y(8) => ALU_OP2_8_port, Y(7) => 
                           ALU_OP2_7_port, Y(6) => ALU_OP2_6_port, Y(5) => 
                           ALU_OP2_5_port, Y(4) => ALU_OP2_4_port, Y(3) => 
                           ALU_OP2_3_port, Y(2) => ALU_OP2_2_port, Y(1) => 
                           ALU_OP2_1_port, Y(0) => ALU_OP2_0_port);
   OUT_MUX : MUX21_GENERIC_NBIT32_2 port map( A(31) => D_DATA_OUT(31), A(30) =>
                           D_DATA_OUT(30), A(29) => D_DATA_OUT(29), A(28) => 
                           D_DATA_OUT(28), A(27) => D_DATA_OUT(27), A(26) => 
                           D_DATA_OUT(26), A(25) => D_DATA_OUT(25), A(24) => 
                           D_DATA_OUT(24), A(23) => D_DATA_OUT(23), A(22) => 
                           D_DATA_OUT(22), A(21) => D_DATA_OUT(21), A(20) => 
                           D_DATA_OUT(20), A(19) => D_DATA_OUT(19), A(18) => 
                           D_DATA_OUT(18), A(17) => D_DATA_OUT(17), A(16) => 
                           D_DATA_OUT(16), A(15) => D_DATA_OUT(15), A(14) => 
                           D_DATA_OUT(14), A(13) => D_DATA_OUT(13), A(12) => 
                           D_DATA_OUT(12), A(11) => D_DATA_OUT(11), A(10) => 
                           D_DATA_OUT(10), A(9) => D_DATA_OUT(9), A(8) => 
                           D_DATA_OUT(8), A(7) => D_DATA_OUT(7), A(6) => 
                           D_DATA_OUT(6), A(5) => D_DATA_OUT(5), A(4) => 
                           D_DATA_OUT(4), A(3) => D_DATA_OUT(3), A(2) => 
                           D_DATA_OUT(2), A(1) => D_DATA_OUT(1), A(0) => 
                           D_DATA_OUT(0), B(31) => current_ALU_OUT2_31_port, 
                           B(30) => current_ALU_OUT2_30_port, B(29) => 
                           current_ALU_OUT2_29_port, B(28) => 
                           current_ALU_OUT2_28_port, B(27) => 
                           current_ALU_OUT2_27_port, B(26) => 
                           current_ALU_OUT2_26_port, B(25) => 
                           current_ALU_OUT2_25_port, B(24) => 
                           current_ALU_OUT2_24_port, B(23) => 
                           current_ALU_OUT2_23_port, B(22) => 
                           current_ALU_OUT2_22_port, B(21) => 
                           current_ALU_OUT2_21_port, B(20) => 
                           current_ALU_OUT2_20_port, B(19) => 
                           current_ALU_OUT2_19_port, B(18) => 
                           current_ALU_OUT2_18_port, B(17) => 
                           current_ALU_OUT2_17_port, B(16) => 
                           current_ALU_OUT2_16_port, B(15) => 
                           current_ALU_OUT2_15_port, B(14) => 
                           current_ALU_OUT2_14_port, B(13) => 
                           current_ALU_OUT2_13_port, B(12) => 
                           current_ALU_OUT2_12_port, B(11) => 
                           current_ALU_OUT2_11_port, B(10) => 
                           current_ALU_OUT2_10_port, B(9) => 
                           current_ALU_OUT2_9_port, B(8) => 
                           current_ALU_OUT2_8_port, B(7) => 
                           current_ALU_OUT2_7_port, B(6) => 
                           current_ALU_OUT2_6_port, B(5) => 
                           current_ALU_OUT2_5_port, B(4) => 
                           current_ALU_OUT2_4_port, B(3) => 
                           current_ALU_OUT2_3_port, B(2) => 
                           current_ALU_OUT2_2_port, B(1) => 
                           current_ALU_OUT2_1_port, B(0) => 
                           current_ALU_OUT2_0_port, SEL => WB_MUX_SEL, Y(31) =>
                           OUT_MUX_DATA_31_port, Y(30) => OUT_MUX_DATA_30_port,
                           Y(29) => OUT_MUX_DATA_29_port, Y(28) => 
                           OUT_MUX_DATA_28_port, Y(27) => OUT_MUX_DATA_27_port,
                           Y(26) => OUT_MUX_DATA_26_port, Y(25) => 
                           OUT_MUX_DATA_25_port, Y(24) => OUT_MUX_DATA_24_port,
                           Y(23) => OUT_MUX_DATA_23_port, Y(22) => 
                           OUT_MUX_DATA_22_port, Y(21) => OUT_MUX_DATA_21_port,
                           Y(20) => OUT_MUX_DATA_20_port, Y(19) => 
                           OUT_MUX_DATA_19_port, Y(18) => OUT_MUX_DATA_18_port,
                           Y(17) => OUT_MUX_DATA_17_port, Y(16) => 
                           OUT_MUX_DATA_16_port, Y(15) => OUT_MUX_DATA_15_port,
                           Y(14) => OUT_MUX_DATA_14_port, Y(13) => 
                           OUT_MUX_DATA_13_port, Y(12) => OUT_MUX_DATA_12_port,
                           Y(11) => OUT_MUX_DATA_11_port, Y(10) => 
                           OUT_MUX_DATA_10_port, Y(9) => OUT_MUX_DATA_9_port, 
                           Y(8) => OUT_MUX_DATA_8_port, Y(7) => 
                           OUT_MUX_DATA_7_port, Y(6) => OUT_MUX_DATA_6_port, 
                           Y(5) => OUT_MUX_DATA_5_port, Y(4) => 
                           OUT_MUX_DATA_4_port, Y(3) => OUT_MUX_DATA_3_port, 
                           Y(2) => OUT_MUX_DATA_2_port, Y(1) => 
                           OUT_MUX_DATA_1_port, Y(0) => OUT_MUX_DATA_0_port);
   JAL_DATA_MUX : MUX21_GENERIC_NBIT32_1 port map( A(31) => 
                           OUT_MUX_DATA_31_port, A(30) => OUT_MUX_DATA_30_port,
                           A(29) => OUT_MUX_DATA_29_port, A(28) => 
                           OUT_MUX_DATA_28_port, A(27) => OUT_MUX_DATA_27_port,
                           A(26) => OUT_MUX_DATA_26_port, A(25) => 
                           OUT_MUX_DATA_25_port, A(24) => OUT_MUX_DATA_24_port,
                           A(23) => OUT_MUX_DATA_23_port, A(22) => 
                           OUT_MUX_DATA_22_port, A(21) => OUT_MUX_DATA_21_port,
                           A(20) => OUT_MUX_DATA_20_port, A(19) => 
                           OUT_MUX_DATA_19_port, A(18) => OUT_MUX_DATA_18_port,
                           A(17) => OUT_MUX_DATA_17_port, A(16) => 
                           OUT_MUX_DATA_16_port, A(15) => OUT_MUX_DATA_15_port,
                           A(14) => OUT_MUX_DATA_14_port, A(13) => 
                           OUT_MUX_DATA_13_port, A(12) => OUT_MUX_DATA_12_port,
                           A(11) => OUT_MUX_DATA_11_port, A(10) => 
                           OUT_MUX_DATA_10_port, A(9) => OUT_MUX_DATA_9_port, 
                           A(8) => OUT_MUX_DATA_8_port, A(7) => 
                           OUT_MUX_DATA_7_port, A(6) => OUT_MUX_DATA_6_port, 
                           A(5) => OUT_MUX_DATA_5_port, A(4) => 
                           OUT_MUX_DATA_4_port, A(3) => OUT_MUX_DATA_3_port, 
                           A(2) => OUT_MUX_DATA_2_port, A(1) => 
                           OUT_MUX_DATA_1_port, A(0) => OUT_MUX_DATA_0_port, 
                           B(31) => current_PC3_31_port, B(30) => 
                           current_PC3_30_port, B(29) => current_PC3_29_port, 
                           B(28) => current_PC3_28_port, B(27) => 
                           current_PC3_27_port, B(26) => current_PC3_26_port, 
                           B(25) => current_PC3_25_port, B(24) => 
                           current_PC3_24_port, B(23) => current_PC3_23_port, 
                           B(22) => current_PC3_22_port, B(21) => 
                           current_PC3_21_port, B(20) => current_PC3_20_port, 
                           B(19) => current_PC3_19_port, B(18) => 
                           current_PC3_18_port, B(17) => current_PC3_17_port, 
                           B(16) => current_PC3_16_port, B(15) => 
                           current_PC3_15_port, B(14) => current_PC3_14_port, 
                           B(13) => current_PC3_13_port, B(12) => 
                           current_PC3_12_port, B(11) => current_PC3_11_port, 
                           B(10) => current_PC3_10_port, B(9) => 
                           current_PC3_9_port, B(8) => current_PC3_8_port, B(7)
                           => current_PC3_7_port, B(6) => current_PC3_6_port, 
                           B(5) => current_PC3_5_port, B(4) => 
                           current_PC3_4_port, B(3) => current_PC3_3_port, B(2)
                           => current_PC3_2_port, B(1) => current_PC3_1_port, 
                           B(0) => current_PC3_0_port, SEL => IS_JAL, Y(31) => 
                           WB_DATA_31_port, Y(30) => WB_DATA_30_port, Y(29) => 
                           WB_DATA_29_port, Y(28) => WB_DATA_28_port, Y(27) => 
                           WB_DATA_27_port, Y(26) => WB_DATA_26_port, Y(25) => 
                           WB_DATA_25_port, Y(24) => WB_DATA_24_port, Y(23) => 
                           WB_DATA_23_port, Y(22) => WB_DATA_22_port, Y(21) => 
                           WB_DATA_21_port, Y(20) => WB_DATA_20_port, Y(19) => 
                           WB_DATA_19_port, Y(18) => WB_DATA_18_port, Y(17) => 
                           WB_DATA_17_port, Y(16) => WB_DATA_16_port, Y(15) => 
                           WB_DATA_15_port, Y(14) => WB_DATA_14_port, Y(13) => 
                           WB_DATA_13_port, Y(12) => WB_DATA_12_port, Y(11) => 
                           WB_DATA_11_port, Y(10) => WB_DATA_10_port, Y(9) => 
                           WB_DATA_9_port, Y(8) => WB_DATA_8_port, Y(7) => 
                           WB_DATA_7_port, Y(6) => WB_DATA_6_port, Y(5) => 
                           WB_DATA_5_port, Y(4) => WB_DATA_4_port, Y(3) => 
                           WB_DATA_3_port, Y(2) => WB_DATA_2_port, Y(1) => 
                           WB_DATA_1_port, Y(0) => WB_DATA_0_port);
   JAL_ADDR_MUX : MUX21_GENERIC_NBIT5_1 port map( A(4) => WB3_OUT_4_port, A(3) 
                           => WB3_OUT_3_port, A(2) => WB3_OUT_2_port, A(1) => 
                           WB3_OUT_1_port, A(0) => WB3_OUT_0_port, B(4) => 
                           X_Logic1_port, B(3) => X_Logic1_port, B(2) => 
                           X_Logic1_port, B(1) => X_Logic1_port, B(0) => 
                           X_Logic1_port, SEL => IS_JAL, Y(4) => WB_ADDR_4_port
                           , Y(3) => WB_ADDR_3_port, Y(2) => WB_ADDR_2_port, 
                           Y(1) => WB_ADDR_1_port, Y(0) => WB_ADDR_0_port);
   PC_ADDER : ADDER_N32 port map( CURR_ADDR(31) => current_PC_31_port, 
                           CURR_ADDR(30) => current_PC_30_port, CURR_ADDR(29) 
                           => current_PC_29_port, CURR_ADDR(28) => 
                           current_PC_28_port, CURR_ADDR(27) => 
                           current_PC_27_port, CURR_ADDR(26) => 
                           current_PC_26_port, CURR_ADDR(25) => 
                           current_PC_25_port, CURR_ADDR(24) => 
                           current_PC_24_port, CURR_ADDR(23) => 
                           current_PC_23_port, CURR_ADDR(22) => 
                           current_PC_22_port, CURR_ADDR(21) => 
                           current_PC_21_port, CURR_ADDR(20) => 
                           current_PC_20_port, CURR_ADDR(19) => 
                           current_PC_19_port, CURR_ADDR(18) => 
                           current_PC_18_port, CURR_ADDR(17) => 
                           current_PC_17_port, CURR_ADDR(16) => 
                           current_PC_16_port, CURR_ADDR(15) => 
                           current_PC_15_port, CURR_ADDR(14) => 
                           current_PC_14_port, CURR_ADDR(13) => 
                           current_PC_13_port, CURR_ADDR(12) => 
                           current_PC_12_port, CURR_ADDR(11) => 
                           current_PC_11_port, CURR_ADDR(10) => 
                           current_PC_10_port, CURR_ADDR(9) => 
                           current_PC_9_port, CURR_ADDR(8) => current_PC_8_port
                           , CURR_ADDR(7) => current_PC_7_port, CURR_ADDR(6) =>
                           current_PC_6_port, CURR_ADDR(5) => current_PC_5_port
                           , CURR_ADDR(4) => current_PC_4_port, CURR_ADDR(3) =>
                           current_PC_3_port, CURR_ADDR(2) => current_PC_2_port
                           , CURR_ADDR(1) => current_PC_1_port, CURR_ADDR(0) =>
                           current_PC_0_port, NEXT_ADDR(31) => next_NPC_31_port
                           , NEXT_ADDR(30) => next_NPC_30_port, NEXT_ADDR(29) 
                           => next_NPC_29_port, NEXT_ADDR(28) => 
                           next_NPC_28_port, NEXT_ADDR(27) => next_NPC_27_port,
                           NEXT_ADDR(26) => next_NPC_26_port, NEXT_ADDR(25) => 
                           next_NPC_25_port, NEXT_ADDR(24) => next_NPC_24_port,
                           NEXT_ADDR(23) => next_NPC_23_port, NEXT_ADDR(22) => 
                           next_NPC_22_port, NEXT_ADDR(21) => next_NPC_21_port,
                           NEXT_ADDR(20) => next_NPC_20_port, NEXT_ADDR(19) => 
                           next_NPC_19_port, NEXT_ADDR(18) => next_NPC_18_port,
                           NEXT_ADDR(17) => next_NPC_17_port, NEXT_ADDR(16) => 
                           next_NPC_16_port, NEXT_ADDR(15) => next_NPC_15_port,
                           NEXT_ADDR(14) => next_NPC_14_port, NEXT_ADDR(13) => 
                           next_NPC_13_port, NEXT_ADDR(12) => next_NPC_12_port,
                           NEXT_ADDR(11) => next_NPC_11_port, NEXT_ADDR(10) => 
                           next_NPC_10_port, NEXT_ADDR(9) => next_NPC_9_port, 
                           NEXT_ADDR(8) => next_NPC_8_port, NEXT_ADDR(7) => 
                           next_NPC_7_port, NEXT_ADDR(6) => next_NPC_6_port, 
                           NEXT_ADDR(5) => next_NPC_5_port, NEXT_ADDR(4) => 
                           next_NPC_4_port, NEXT_ADDR(3) => next_NPC_3_port, 
                           NEXT_ADDR(2) => next_NPC_2_port, NEXT_ADDR(1) => 
                           next_NPC_1_port, NEXT_ADDR(0) => next_NPC_0_port);
   RF : REGISTER_FILE_NBIT32_NREG32 port map( CLK => CLK, RST => RST, EN => 
                           X_Logic1_port, RD1 => RegA_LATCH_EN, RD2 => 
                           RegB_LATCH_EN, WR => RF_WE, ADD_WR(4) => 
                           WB_ADDR_4_port, ADD_WR(3) => WB_ADDR_3_port, 
                           ADD_WR(2) => WB_ADDR_2_port, ADD_WR(1) => 
                           WB_ADDR_1_port, ADD_WR(0) => WB_ADDR_0_port, 
                           ADD_RD1(4) => current_IW_25_port, ADD_RD1(3) => 
                           current_IW_24_port, ADD_RD1(2) => current_IW_23_port
                           , ADD_RD1(1) => current_IW_22_port, ADD_RD1(0) => 
                           current_IW_21_port, ADD_RD2(4) => current_IW_20_port
                           , ADD_RD2(3) => current_IW_19_port, ADD_RD2(2) => 
                           current_IW_18_port, ADD_RD2(1) => current_IW_17_port
                           , ADD_RD2(0) => current_IW_16_port, DATAIN(31) => 
                           WB_DATA_31_port, DATAIN(30) => WB_DATA_30_port, 
                           DATAIN(29) => WB_DATA_29_port, DATAIN(28) => 
                           WB_DATA_28_port, DATAIN(27) => WB_DATA_27_port, 
                           DATAIN(26) => WB_DATA_26_port, DATAIN(25) => 
                           WB_DATA_25_port, DATAIN(24) => WB_DATA_24_port, 
                           DATAIN(23) => WB_DATA_23_port, DATAIN(22) => 
                           WB_DATA_22_port, DATAIN(21) => WB_DATA_21_port, 
                           DATAIN(20) => WB_DATA_20_port, DATAIN(19) => 
                           WB_DATA_19_port, DATAIN(18) => WB_DATA_18_port, 
                           DATAIN(17) => WB_DATA_17_port, DATAIN(16) => 
                           WB_DATA_16_port, DATAIN(15) => WB_DATA_15_port, 
                           DATAIN(14) => WB_DATA_14_port, DATAIN(13) => 
                           WB_DATA_13_port, DATAIN(12) => WB_DATA_12_port, 
                           DATAIN(11) => WB_DATA_11_port, DATAIN(10) => 
                           WB_DATA_10_port, DATAIN(9) => WB_DATA_9_port, 
                           DATAIN(8) => WB_DATA_8_port, DATAIN(7) => 
                           WB_DATA_7_port, DATAIN(6) => WB_DATA_6_port, 
                           DATAIN(5) => WB_DATA_5_port, DATAIN(4) => 
                           WB_DATA_4_port, DATAIN(3) => WB_DATA_3_port, 
                           DATAIN(2) => WB_DATA_2_port, DATAIN(1) => 
                           WB_DATA_1_port, DATAIN(0) => WB_DATA_0_port, 
                           OUT1(31) => A_OUT_31_port, OUT1(30) => A_OUT_30_port
                           , OUT1(29) => A_OUT_29_port, OUT1(28) => 
                           A_OUT_28_port, OUT1(27) => A_OUT_27_port, OUT1(26) 
                           => A_OUT_26_port, OUT1(25) => A_OUT_25_port, 
                           OUT1(24) => A_OUT_24_port, OUT1(23) => A_OUT_23_port
                           , OUT1(22) => A_OUT_22_port, OUT1(21) => 
                           A_OUT_21_port, OUT1(20) => A_OUT_20_port, OUT1(19) 
                           => A_OUT_19_port, OUT1(18) => A_OUT_18_port, 
                           OUT1(17) => A_OUT_17_port, OUT1(16) => A_OUT_16_port
                           , OUT1(15) => A_OUT_15_port, OUT1(14) => 
                           A_OUT_14_port, OUT1(13) => A_OUT_13_port, OUT1(12) 
                           => A_OUT_12_port, OUT1(11) => A_OUT_11_port, 
                           OUT1(10) => A_OUT_10_port, OUT1(9) => A_OUT_9_port, 
                           OUT1(8) => A_OUT_8_port, OUT1(7) => A_OUT_7_port, 
                           OUT1(6) => A_OUT_6_port, OUT1(5) => A_OUT_5_port, 
                           OUT1(4) => A_OUT_4_port, OUT1(3) => A_OUT_3_port, 
                           OUT1(2) => A_OUT_2_port, OUT1(1) => A_OUT_1_port, 
                           OUT1(0) => A_OUT_0_port, OUT2(31) => B_OUT_31_port, 
                           OUT2(30) => B_OUT_30_port, OUT2(29) => B_OUT_29_port
                           , OUT2(28) => B_OUT_28_port, OUT2(27) => 
                           B_OUT_27_port, OUT2(26) => B_OUT_26_port, OUT2(25) 
                           => B_OUT_25_port, OUT2(24) => B_OUT_24_port, 
                           OUT2(23) => B_OUT_23_port, OUT2(22) => B_OUT_22_port
                           , OUT2(21) => B_OUT_21_port, OUT2(20) => 
                           B_OUT_20_port, OUT2(19) => B_OUT_19_port, OUT2(18) 
                           => B_OUT_18_port, OUT2(17) => B_OUT_17_port, 
                           OUT2(16) => B_OUT_16_port, OUT2(15) => B_OUT_15_port
                           , OUT2(14) => B_OUT_14_port, OUT2(13) => 
                           B_OUT_13_port, OUT2(12) => B_OUT_12_port, OUT2(11) 
                           => B_OUT_11_port, OUT2(10) => B_OUT_10_port, OUT2(9)
                           => B_OUT_9_port, OUT2(8) => B_OUT_8_port, OUT2(7) =>
                           B_OUT_7_port, OUT2(6) => B_OUT_6_port, OUT2(5) => 
                           B_OUT_5_port, OUT2(4) => B_OUT_4_port, OUT2(3) => 
                           B_OUT_3_port, OUT2(2) => B_OUT_2_port, OUT2(1) => 
                           B_OUT_1_port, OUT2(0) => B_OUT_0_port);
   EXT : EXTENDER_NBIT32_IMM_MIN16_IMM_MAX26 port map( NOT_EXT_IMM(25) => 
                           IMM_IN_25_port, NOT_EXT_IMM(24) => IMM_IN_24_port, 
                           NOT_EXT_IMM(23) => IMM_IN_23_port, NOT_EXT_IMM(22) 
                           => IMM_IN_22_port, NOT_EXT_IMM(21) => IMM_IN_21_port
                           , NOT_EXT_IMM(20) => IMM_IN_20_port, NOT_EXT_IMM(19)
                           => IMM_IN_19_port, NOT_EXT_IMM(18) => IMM_IN_18_port
                           , NOT_EXT_IMM(17) => IMM_IN_17_port, NOT_EXT_IMM(16)
                           => IMM_IN_16_port, NOT_EXT_IMM(15) => IMM_IN_15_port
                           , NOT_EXT_IMM(14) => IMM_IN_14_port, NOT_EXT_IMM(13)
                           => IMM_IN_13_port, NOT_EXT_IMM(12) => IMM_IN_12_port
                           , NOT_EXT_IMM(11) => IMM_IN_11_port, NOT_EXT_IMM(10)
                           => IMM_IN_10_port, NOT_EXT_IMM(9) => IMM_IN_9_port, 
                           NOT_EXT_IMM(8) => IMM_IN_8_port, NOT_EXT_IMM(7) => 
                           IMM_IN_7_port, NOT_EXT_IMM(6) => IMM_IN_6_port, 
                           NOT_EXT_IMM(5) => IMM_IN_5_port, NOT_EXT_IMM(4) => 
                           IMM_IN_4_port, NOT_EXT_IMM(3) => IMM_IN_3_port, 
                           NOT_EXT_IMM(2) => IMM_IN_2_port, NOT_EXT_IMM(1) => 
                           IMM_IN_1_port, NOT_EXT_IMM(0) => IMM_IN_0_port, 
                           SIGNED_IMM => SIGNED_IMM, IS_JUMP => IS_JUMP, 
                           EXT_IMM(31) => IMM_OUT_31_port, EXT_IMM(30) => 
                           IMM_OUT_30_port, EXT_IMM(29) => IMM_OUT_29_port, 
                           EXT_IMM(28) => IMM_OUT_28_port, EXT_IMM(27) => 
                           IMM_OUT_27_port, EXT_IMM(26) => IMM_OUT_26_port, 
                           EXT_IMM(25) => IMM_OUT_25_port, EXT_IMM(24) => 
                           IMM_OUT_24_port, EXT_IMM(23) => IMM_OUT_23_port, 
                           EXT_IMM(22) => IMM_OUT_22_port, EXT_IMM(21) => 
                           IMM_OUT_21_port, EXT_IMM(20) => IMM_OUT_20_port, 
                           EXT_IMM(19) => IMM_OUT_19_port, EXT_IMM(18) => 
                           IMM_OUT_18_port, EXT_IMM(17) => IMM_OUT_17_port, 
                           EXT_IMM(16) => IMM_OUT_16_port, EXT_IMM(15) => 
                           IMM_OUT_15_port, EXT_IMM(14) => IMM_OUT_14_port, 
                           EXT_IMM(13) => IMM_OUT_13_port, EXT_IMM(12) => 
                           IMM_OUT_12_port, EXT_IMM(11) => IMM_OUT_11_port, 
                           EXT_IMM(10) => IMM_OUT_10_port, EXT_IMM(9) => 
                           IMM_OUT_9_port, EXT_IMM(8) => IMM_OUT_8_port, 
                           EXT_IMM(7) => IMM_OUT_7_port, EXT_IMM(6) => 
                           IMM_OUT_6_port, EXT_IMM(5) => IMM_OUT_5_port, 
                           EXT_IMM(4) => IMM_OUT_4_port, EXT_IMM(3) => 
                           IMM_OUT_3_port, EXT_IMM(2) => IMM_OUT_2_port, 
                           EXT_IMM(1) => IMM_OUT_1_port, EXT_IMM(0) => 
                           IMM_OUT_0_port);
   ALU_i : ALU_N32 port map( FUNC(0) => ALU_OPCODE(0), FUNC(1) => ALU_OPCODE(1)
                           , FUNC(2) => ALU_OPCODE(2), FUNC(3) => ALU_OPCODE(3)
                           , DATA1(31) => ALU_OP1_31_port, DATA1(30) => 
                           ALU_OP1_30_port, DATA1(29) => ALU_OP1_29_port, 
                           DATA1(28) => ALU_OP1_28_port, DATA1(27) => 
                           ALU_OP1_27_port, DATA1(26) => ALU_OP1_26_port, 
                           DATA1(25) => ALU_OP1_25_port, DATA1(24) => 
                           ALU_OP1_24_port, DATA1(23) => ALU_OP1_23_port, 
                           DATA1(22) => ALU_OP1_22_port, DATA1(21) => 
                           ALU_OP1_21_port, DATA1(20) => ALU_OP1_20_port, 
                           DATA1(19) => ALU_OP1_19_port, DATA1(18) => 
                           ALU_OP1_18_port, DATA1(17) => ALU_OP1_17_port, 
                           DATA1(16) => ALU_OP1_16_port, DATA1(15) => 
                           ALU_OP1_15_port, DATA1(14) => ALU_OP1_14_port, 
                           DATA1(13) => ALU_OP1_13_port, DATA1(12) => 
                           ALU_OP1_12_port, DATA1(11) => ALU_OP1_11_port, 
                           DATA1(10) => ALU_OP1_10_port, DATA1(9) => 
                           ALU_OP1_9_port, DATA1(8) => ALU_OP1_8_port, DATA1(7)
                           => ALU_OP1_7_port, DATA1(6) => ALU_OP1_6_port, 
                           DATA1(5) => ALU_OP1_5_port, DATA1(4) => 
                           ALU_OP1_4_port, DATA1(3) => ALU_OP1_3_port, DATA1(2)
                           => ALU_OP1_2_port, DATA1(1) => ALU_OP1_1_port, 
                           DATA1(0) => ALU_OP1_0_port, DATA2(31) => 
                           ALU_OP2_31_port, DATA2(30) => ALU_OP2_30_port, 
                           DATA2(29) => ALU_OP2_29_port, DATA2(28) => 
                           ALU_OP2_28_port, DATA2(27) => ALU_OP2_27_port, 
                           DATA2(26) => ALU_OP2_26_port, DATA2(25) => 
                           ALU_OP2_25_port, DATA2(24) => ALU_OP2_24_port, 
                           DATA2(23) => ALU_OP2_23_port, DATA2(22) => 
                           ALU_OP2_22_port, DATA2(21) => ALU_OP2_21_port, 
                           DATA2(20) => ALU_OP2_20_port, DATA2(19) => 
                           ALU_OP2_19_port, DATA2(18) => ALU_OP2_18_port, 
                           DATA2(17) => ALU_OP2_17_port, DATA2(16) => 
                           ALU_OP2_16_port, DATA2(15) => ALU_OP2_15_port, 
                           DATA2(14) => ALU_OP2_14_port, DATA2(13) => 
                           ALU_OP2_13_port, DATA2(12) => ALU_OP2_12_port, 
                           DATA2(11) => ALU_OP2_11_port, DATA2(10) => 
                           ALU_OP2_10_port, DATA2(9) => ALU_OP2_9_port, 
                           DATA2(8) => ALU_OP2_8_port, DATA2(7) => 
                           ALU_OP2_7_port, DATA2(6) => ALU_OP2_6_port, DATA2(5)
                           => ALU_OP2_5_port, DATA2(4) => ALU_OP2_4_port, 
                           DATA2(3) => ALU_OP2_3_port, DATA2(2) => 
                           ALU_OP2_2_port, DATA2(1) => ALU_OP2_1_port, DATA2(0)
                           => ALU_OP2_0_port, OUTALU(31) => 
                           next_ALU_OUT_31_port, OUTALU(30) => 
                           next_ALU_OUT_30_port, OUTALU(29) => 
                           next_ALU_OUT_29_port, OUTALU(28) => 
                           next_ALU_OUT_28_port, OUTALU(27) => 
                           next_ALU_OUT_27_port, OUTALU(26) => 
                           next_ALU_OUT_26_port, OUTALU(25) => 
                           next_ALU_OUT_25_port, OUTALU(24) => 
                           next_ALU_OUT_24_port, OUTALU(23) => 
                           next_ALU_OUT_23_port, OUTALU(22) => 
                           next_ALU_OUT_22_port, OUTALU(21) => 
                           next_ALU_OUT_21_port, OUTALU(20) => 
                           next_ALU_OUT_20_port, OUTALU(19) => 
                           next_ALU_OUT_19_port, OUTALU(18) => 
                           next_ALU_OUT_18_port, OUTALU(17) => 
                           next_ALU_OUT_17_port, OUTALU(16) => 
                           next_ALU_OUT_16_port, OUTALU(15) => 
                           next_ALU_OUT_15_port, OUTALU(14) => 
                           next_ALU_OUT_14_port, OUTALU(13) => 
                           next_ALU_OUT_13_port, OUTALU(12) => 
                           next_ALU_OUT_12_port, OUTALU(11) => 
                           next_ALU_OUT_11_port, OUTALU(10) => 
                           next_ALU_OUT_10_port, OUTALU(9) => 
                           next_ALU_OUT_9_port, OUTALU(8) => 
                           next_ALU_OUT_8_port, OUTALU(7) => 
                           next_ALU_OUT_7_port, OUTALU(6) => 
                           next_ALU_OUT_6_port, OUTALU(5) => 
                           next_ALU_OUT_5_port, OUTALU(4) => 
                           next_ALU_OUT_4_port, OUTALU(3) => 
                           next_ALU_OUT_3_port, OUTALU(2) => 
                           next_ALU_OUT_2_port, OUTALU(1) => 
                           next_ALU_OUT_1_port, OUTALU(0) => 
                           next_ALU_OUT_0_port);
   U3 : AND2_X1 port map( A1 => PC_LATCH_EN, A2 => PC_BUS_9_port, ZN => 
                           current_PC_9_port);
   U4 : AND2_X1 port map( A1 => PC_BUS_8_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_8_port);
   U5 : AND2_X1 port map( A1 => PC_BUS_7_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_7_port);
   U6 : AND2_X1 port map( A1 => PC_BUS_6_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_6_port);
   U7 : AND2_X1 port map( A1 => PC_BUS_5_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_5_port);
   U8 : AND2_X1 port map( A1 => PC_BUS_4_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_4_port);
   U9 : AND2_X1 port map( A1 => PC_BUS_3_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_3_port);
   U10 : AND2_X1 port map( A1 => PC_BUS_31_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_31_port);
   U11 : AND2_X1 port map( A1 => PC_BUS_30_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_30_port);
   U12 : AND2_X1 port map( A1 => PC_BUS_2_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_2_port);
   U13 : AND2_X1 port map( A1 => PC_BUS_29_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_29_port);
   U14 : AND2_X1 port map( A1 => PC_BUS_28_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_28_port);
   U15 : AND2_X1 port map( A1 => PC_BUS_27_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_27_port);
   U16 : AND2_X1 port map( A1 => PC_BUS_26_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_26_port);
   U17 : AND2_X1 port map( A1 => PC_BUS_25_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_25_port);
   U18 : AND2_X1 port map( A1 => PC_BUS_24_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_24_port);
   U19 : AND2_X1 port map( A1 => PC_BUS_23_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_23_port);
   U20 : AND2_X1 port map( A1 => PC_BUS_22_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_22_port);
   U21 : AND2_X1 port map( A1 => PC_BUS_21_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_21_port);
   U22 : AND2_X1 port map( A1 => PC_BUS_20_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_20_port);
   U23 : AND2_X1 port map( A1 => PC_BUS_1_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_1_port);
   U24 : AND2_X1 port map( A1 => PC_BUS_19_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_19_port);
   U25 : AND2_X1 port map( A1 => PC_BUS_18_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_18_port);
   U26 : AND2_X1 port map( A1 => PC_BUS_17_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_17_port);
   U27 : AND2_X1 port map( A1 => PC_BUS_16_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_16_port);
   U28 : AND2_X1 port map( A1 => PC_BUS_15_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_15_port);
   U29 : AND2_X1 port map( A1 => PC_BUS_14_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_14_port);
   U30 : AND2_X1 port map( A1 => PC_BUS_13_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_13_port);
   U31 : AND2_X1 port map( A1 => PC_BUS_12_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_12_port);
   U32 : AND2_X1 port map( A1 => PC_BUS_11_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_11_port);
   U33 : AND2_X1 port map( A1 => PC_BUS_10_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_10_port);
   U34 : AND2_X1 port map( A1 => PC_BUS_0_port, A2 => PC_LATCH_EN, ZN => 
                           current_PC_0_port);

end SYN_STRUCTURE;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REG_GENERIC_NBIT32_0 is

   port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 downto
         0);  DATA_OUT : out std_logic_vector (31 downto 0));

end REG_GENERIC_NBIT32_0;

architecture SYN_BEHAVIOR of REG_GENERIC_NBIT32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   DATA_OUT_reg_31_inst : DFF_X1 port map( D => n68, CK => CLK, Q => 
                           DATA_OUT(31), QN => n67);
   DATA_OUT_reg_30_inst : DFF_X1 port map( D => n69, CK => CLK, Q => 
                           DATA_OUT(30), QN => n66);
   DATA_OUT_reg_29_inst : DFF_X1 port map( D => n70, CK => CLK, Q => 
                           DATA_OUT(29), QN => n65);
   DATA_OUT_reg_28_inst : DFF_X1 port map( D => n71, CK => CLK, Q => 
                           DATA_OUT(28), QN => n64);
   DATA_OUT_reg_27_inst : DFF_X1 port map( D => n72, CK => CLK, Q => 
                           DATA_OUT(27), QN => n63);
   DATA_OUT_reg_26_inst : DFF_X1 port map( D => n73, CK => CLK, Q => 
                           DATA_OUT(26), QN => n62);
   DATA_OUT_reg_25_inst : DFF_X1 port map( D => n74, CK => CLK, Q => 
                           DATA_OUT(25), QN => n61);
   DATA_OUT_reg_24_inst : DFF_X1 port map( D => n75, CK => CLK, Q => 
                           DATA_OUT(24), QN => n60);
   DATA_OUT_reg_23_inst : DFF_X1 port map( D => n76, CK => CLK, Q => 
                           DATA_OUT(23), QN => n59);
   DATA_OUT_reg_22_inst : DFF_X1 port map( D => n77, CK => CLK, Q => 
                           DATA_OUT(22), QN => n58);
   DATA_OUT_reg_21_inst : DFF_X1 port map( D => n78, CK => CLK, Q => 
                           DATA_OUT(21), QN => n57);
   DATA_OUT_reg_20_inst : DFF_X1 port map( D => n79, CK => CLK, Q => 
                           DATA_OUT(20), QN => n56);
   DATA_OUT_reg_19_inst : DFF_X1 port map( D => n80, CK => CLK, Q => 
                           DATA_OUT(19), QN => n55);
   DATA_OUT_reg_18_inst : DFF_X1 port map( D => n81, CK => CLK, Q => 
                           DATA_OUT(18), QN => n54);
   DATA_OUT_reg_17_inst : DFF_X1 port map( D => n82, CK => CLK, Q => 
                           DATA_OUT(17), QN => n53);
   DATA_OUT_reg_16_inst : DFF_X1 port map( D => n83, CK => CLK, Q => 
                           DATA_OUT(16), QN => n52);
   DATA_OUT_reg_15_inst : DFF_X1 port map( D => n84, CK => CLK, Q => 
                           DATA_OUT(15), QN => n51);
   DATA_OUT_reg_14_inst : DFF_X1 port map( D => n85, CK => CLK, Q => 
                           DATA_OUT(14), QN => n50);
   DATA_OUT_reg_13_inst : DFF_X1 port map( D => n86, CK => CLK, Q => 
                           DATA_OUT(13), QN => n49);
   DATA_OUT_reg_12_inst : DFF_X1 port map( D => n87, CK => CLK, Q => 
                           DATA_OUT(12), QN => n48);
   DATA_OUT_reg_11_inst : DFF_X1 port map( D => n88, CK => CLK, Q => 
                           DATA_OUT(11), QN => n47);
   DATA_OUT_reg_10_inst : DFF_X1 port map( D => n89, CK => CLK, Q => 
                           DATA_OUT(10), QN => n46);
   DATA_OUT_reg_9_inst : DFF_X1 port map( D => n90, CK => CLK, Q => DATA_OUT(9)
                           , QN => n45);
   DATA_OUT_reg_8_inst : DFF_X1 port map( D => n91, CK => CLK, Q => DATA_OUT(8)
                           , QN => n44);
   DATA_OUT_reg_7_inst : DFF_X1 port map( D => n92, CK => CLK, Q => DATA_OUT(7)
                           , QN => n43);
   DATA_OUT_reg_6_inst : DFF_X1 port map( D => n93, CK => CLK, Q => DATA_OUT(6)
                           , QN => n42);
   DATA_OUT_reg_5_inst : DFF_X1 port map( D => n94, CK => CLK, Q => DATA_OUT(5)
                           , QN => n41);
   DATA_OUT_reg_4_inst : DFF_X1 port map( D => n95, CK => CLK, Q => DATA_OUT(4)
                           , QN => n40);
   DATA_OUT_reg_3_inst : DFF_X1 port map( D => n96, CK => CLK, Q => DATA_OUT(3)
                           , QN => n39);
   DATA_OUT_reg_2_inst : DFF_X1 port map( D => n97, CK => CLK, Q => DATA_OUT(2)
                           , QN => n38);
   DATA_OUT_reg_1_inst : DFF_X1 port map( D => n98, CK => CLK, Q => DATA_OUT(1)
                           , QN => n37);
   DATA_OUT_reg_0_inst : DFF_X1 port map( D => n99, CK => CLK, Q => DATA_OUT(0)
                           , QN => n36);
   U3 : NAND2_X2 port map( A1 => RST, A2 => n1, ZN => n2);
   U4 : NAND2_X2 port map( A1 => n35, A2 => RST, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => DATA_IN(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => DATA_IN(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => DATA_IN(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => DATA_IN(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => DATA_IN(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => DATA_IN(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => DATA_IN(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => DATA_IN(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => DATA_IN(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => DATA_IN(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => DATA_IN(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => DATA_IN(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => DATA_IN(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => DATA_IN(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => DATA_IN(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => DATA_IN(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => DATA_IN(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => DATA_IN(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => DATA_IN(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => DATA_IN(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => DATA_IN(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => DATA_IN(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => DATA_IN(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => DATA_IN(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => DATA_IN(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => DATA_IN(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => DATA_IN(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => DATA_IN(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => DATA_IN(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => DATA_IN(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => DATA_IN(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => DATA_IN(0), ZN => n34);
   U69 : INV_X1 port map( A => EN, ZN => n35);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( CLK, RST : in std_logic;  I_ADDR : out std_logic_vector (31 downto 0);
         I_DATA : in std_logic_vector (31 downto 0);  D_RR, D_WR : out 
         std_logic;  D_ADDR : out std_logic_vector (5 downto 0);  D_DATA_IN : 
         out std_logic_vector (31 downto 0);  D_DATA_OUT : in std_logic_vector 
         (31 downto 0));

end DLX;

architecture SYN_DLX_RTL of DLX is

   component dlx_cu
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
            EQ_COND, IS_JUMP : out std_logic;  ALU_OPCODE : out 
            std_logic_vector (0 to 3);  DRAM_WE, LMD_LATCH_EN, JUMP_EN, 
            PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE : out std_logic);
   end component;
   
   component DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64
      port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
            EQ_COND, IS_JUMP : in std_logic;  ALU_OPCODE : in std_logic_vector 
            (0 to 3);  JUMP_EN, PC_LATCH_EN, IS_JAL, WB_MUX_SEL, RF_WE : in 
            std_logic;  D_ADDR : out std_logic_vector (5 downto 0);  D_DATA_IN 
            : out std_logic_vector (31 downto 0);  D_DATA_OUT, PC_IN : in 
            std_logic_vector (31 downto 0);  PC_BUS : out std_logic_vector (31 
            downto 0));
   end component;
   
   component REG_GENERIC_NBIT32_0
      port( CLK, RST, EN : in std_logic;  DATA_IN : in std_logic_vector (31 
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal I_ADDR_31_port, I_ADDR_30_port, I_ADDR_29_port, I_ADDR_28_port, 
      I_ADDR_27_port, I_ADDR_26_port, I_ADDR_25_port, I_ADDR_24_port, 
      I_ADDR_23_port, I_ADDR_22_port, I_ADDR_21_port, I_ADDR_20_port, 
      I_ADDR_19_port, I_ADDR_18_port, I_ADDR_17_port, I_ADDR_16_port, 
      I_ADDR_15_port, I_ADDR_14_port, I_ADDR_13_port, I_ADDR_12_port, 
      I_ADDR_11_port, I_ADDR_10_port, I_ADDR_9_port, I_ADDR_8_port, 
      I_ADDR_7_port, I_ADDR_6_port, I_ADDR_5_port, I_ADDR_4_port, I_ADDR_3_port
      , I_ADDR_2_port, I_ADDR_1_port, I_ADDR_0_port, PC_LATCH_EN, 
      PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, IR_LATCH_EN, NPC_LATCH_EN,
      RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, SIGNED_IMM, MUXA_SEL, 
      MUXB_SEL, ALU_OUTREG_EN, EQ_COND, IS_JUMP, ALU_OPCODE_3_port, 
      ALU_OPCODE_2_port, ALU_OPCODE_1_port, ALU_OPCODE_0_port, JUMP_EN, IS_JAL,
      WB_MUX_SEL, RF_WE : std_logic;

begin
   I_ADDR <= ( I_ADDR_31_port, I_ADDR_30_port, I_ADDR_29_port, I_ADDR_28_port, 
      I_ADDR_27_port, I_ADDR_26_port, I_ADDR_25_port, I_ADDR_24_port, 
      I_ADDR_23_port, I_ADDR_22_port, I_ADDR_21_port, I_ADDR_20_port, 
      I_ADDR_19_port, I_ADDR_18_port, I_ADDR_17_port, I_ADDR_16_port, 
      I_ADDR_15_port, I_ADDR_14_port, I_ADDR_13_port, I_ADDR_12_port, 
      I_ADDR_11_port, I_ADDR_10_port, I_ADDR_9_port, I_ADDR_8_port, 
      I_ADDR_7_port, I_ADDR_6_port, I_ADDR_5_port, I_ADDR_4_port, I_ADDR_3_port
      , I_ADDR_2_port, I_ADDR_1_port, I_ADDR_0_port );
   
   PC_REG : REG_GENERIC_NBIT32_0 port map( CLK => CLK, RST => RST, EN => 
                           PC_LATCH_EN, DATA_IN(31) => PC_BUS_31_port, 
                           DATA_IN(30) => PC_BUS_30_port, DATA_IN(29) => 
                           PC_BUS_29_port, DATA_IN(28) => PC_BUS_28_port, 
                           DATA_IN(27) => PC_BUS_27_port, DATA_IN(26) => 
                           PC_BUS_26_port, DATA_IN(25) => PC_BUS_25_port, 
                           DATA_IN(24) => PC_BUS_24_port, DATA_IN(23) => 
                           PC_BUS_23_port, DATA_IN(22) => PC_BUS_22_port, 
                           DATA_IN(21) => PC_BUS_21_port, DATA_IN(20) => 
                           PC_BUS_20_port, DATA_IN(19) => PC_BUS_19_port, 
                           DATA_IN(18) => PC_BUS_18_port, DATA_IN(17) => 
                           PC_BUS_17_port, DATA_IN(16) => PC_BUS_16_port, 
                           DATA_IN(15) => PC_BUS_15_port, DATA_IN(14) => 
                           PC_BUS_14_port, DATA_IN(13) => PC_BUS_13_port, 
                           DATA_IN(12) => PC_BUS_12_port, DATA_IN(11) => 
                           PC_BUS_11_port, DATA_IN(10) => PC_BUS_10_port, 
                           DATA_IN(9) => PC_BUS_9_port, DATA_IN(8) => 
                           PC_BUS_8_port, DATA_IN(7) => PC_BUS_7_port, 
                           DATA_IN(6) => PC_BUS_6_port, DATA_IN(5) => 
                           PC_BUS_5_port, DATA_IN(4) => PC_BUS_4_port, 
                           DATA_IN(3) => PC_BUS_3_port, DATA_IN(2) => 
                           PC_BUS_2_port, DATA_IN(1) => PC_BUS_1_port, 
                           DATA_IN(0) => PC_BUS_0_port, DATA_OUT(31) => 
                           I_ADDR_31_port, DATA_OUT(30) => I_ADDR_30_port, 
                           DATA_OUT(29) => I_ADDR_29_port, DATA_OUT(28) => 
                           I_ADDR_28_port, DATA_OUT(27) => I_ADDR_27_port, 
                           DATA_OUT(26) => I_ADDR_26_port, DATA_OUT(25) => 
                           I_ADDR_25_port, DATA_OUT(24) => I_ADDR_24_port, 
                           DATA_OUT(23) => I_ADDR_23_port, DATA_OUT(22) => 
                           I_ADDR_22_port, DATA_OUT(21) => I_ADDR_21_port, 
                           DATA_OUT(20) => I_ADDR_20_port, DATA_OUT(19) => 
                           I_ADDR_19_port, DATA_OUT(18) => I_ADDR_18_port, 
                           DATA_OUT(17) => I_ADDR_17_port, DATA_OUT(16) => 
                           I_ADDR_16_port, DATA_OUT(15) => I_ADDR_15_port, 
                           DATA_OUT(14) => I_ADDR_14_port, DATA_OUT(13) => 
                           I_ADDR_13_port, DATA_OUT(12) => I_ADDR_12_port, 
                           DATA_OUT(11) => I_ADDR_11_port, DATA_OUT(10) => 
                           I_ADDR_10_port, DATA_OUT(9) => I_ADDR_9_port, 
                           DATA_OUT(8) => I_ADDR_8_port, DATA_OUT(7) => 
                           I_ADDR_7_port, DATA_OUT(6) => I_ADDR_6_port, 
                           DATA_OUT(5) => I_ADDR_5_port, DATA_OUT(4) => 
                           I_ADDR_4_port, DATA_OUT(3) => I_ADDR_3_port, 
                           DATA_OUT(2) => I_ADDR_2_port, DATA_OUT(1) => 
                           I_ADDR_1_port, DATA_OUT(0) => I_ADDR_0_port);
   DP : DataPath_BASIC_N32_IR_SIZE32_RF_SIZE32_DRAM_SIZE64 port map( CLK => CLK
                           , RST => RST, IR_IN(31) => I_DATA(31), IR_IN(30) => 
                           I_DATA(30), IR_IN(29) => I_DATA(29), IR_IN(28) => 
                           I_DATA(28), IR_IN(27) => I_DATA(27), IR_IN(26) => 
                           I_DATA(26), IR_IN(25) => I_DATA(25), IR_IN(24) => 
                           I_DATA(24), IR_IN(23) => I_DATA(23), IR_IN(22) => 
                           I_DATA(22), IR_IN(21) => I_DATA(21), IR_IN(20) => 
                           I_DATA(20), IR_IN(19) => I_DATA(19), IR_IN(18) => 
                           I_DATA(18), IR_IN(17) => I_DATA(17), IR_IN(16) => 
                           I_DATA(16), IR_IN(15) => I_DATA(15), IR_IN(14) => 
                           I_DATA(14), IR_IN(13) => I_DATA(13), IR_IN(12) => 
                           I_DATA(12), IR_IN(11) => I_DATA(11), IR_IN(10) => 
                           I_DATA(10), IR_IN(9) => I_DATA(9), IR_IN(8) => 
                           I_DATA(8), IR_IN(7) => I_DATA(7), IR_IN(6) => 
                           I_DATA(6), IR_IN(5) => I_DATA(5), IR_IN(4) => 
                           I_DATA(4), IR_IN(3) => I_DATA(3), IR_IN(2) => 
                           I_DATA(2), IR_IN(1) => I_DATA(1), IR_IN(0) => 
                           I_DATA(0), IR_LATCH_EN => IR_LATCH_EN, NPC_LATCH_EN 
                           => NPC_LATCH_EN, RegA_LATCH_EN => RegA_LATCH_EN, 
                           RegB_LATCH_EN => RegB_LATCH_EN, RegIMM_LATCH_EN => 
                           RegIMM_LATCH_EN, SIGNED_IMM => SIGNED_IMM, MUXA_SEL 
                           => MUXA_SEL, MUXB_SEL => MUXB_SEL, ALU_OUTREG_EN => 
                           ALU_OUTREG_EN, EQ_COND => EQ_COND, IS_JUMP => 
                           IS_JUMP, ALU_OPCODE(0) => ALU_OPCODE_3_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_2_port, ALU_OPCODE(2) =>
                           ALU_OPCODE_1_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_0_port, JUMP_EN => JUMP_EN, PC_LATCH_EN 
                           => PC_LATCH_EN, IS_JAL => IS_JAL, WB_MUX_SEL => 
                           WB_MUX_SEL, RF_WE => RF_WE, D_ADDR(5) => D_ADDR(5), 
                           D_ADDR(4) => D_ADDR(4), D_ADDR(3) => D_ADDR(3), 
                           D_ADDR(2) => D_ADDR(2), D_ADDR(1) => D_ADDR(1), 
                           D_ADDR(0) => D_ADDR(0), D_DATA_IN(31) => 
                           D_DATA_IN(31), D_DATA_IN(30) => D_DATA_IN(30), 
                           D_DATA_IN(29) => D_DATA_IN(29), D_DATA_IN(28) => 
                           D_DATA_IN(28), D_DATA_IN(27) => D_DATA_IN(27), 
                           D_DATA_IN(26) => D_DATA_IN(26), D_DATA_IN(25) => 
                           D_DATA_IN(25), D_DATA_IN(24) => D_DATA_IN(24), 
                           D_DATA_IN(23) => D_DATA_IN(23), D_DATA_IN(22) => 
                           D_DATA_IN(22), D_DATA_IN(21) => D_DATA_IN(21), 
                           D_DATA_IN(20) => D_DATA_IN(20), D_DATA_IN(19) => 
                           D_DATA_IN(19), D_DATA_IN(18) => D_DATA_IN(18), 
                           D_DATA_IN(17) => D_DATA_IN(17), D_DATA_IN(16) => 
                           D_DATA_IN(16), D_DATA_IN(15) => D_DATA_IN(15), 
                           D_DATA_IN(14) => D_DATA_IN(14), D_DATA_IN(13) => 
                           D_DATA_IN(13), D_DATA_IN(12) => D_DATA_IN(12), 
                           D_DATA_IN(11) => D_DATA_IN(11), D_DATA_IN(10) => 
                           D_DATA_IN(10), D_DATA_IN(9) => D_DATA_IN(9), 
                           D_DATA_IN(8) => D_DATA_IN(8), D_DATA_IN(7) => 
                           D_DATA_IN(7), D_DATA_IN(6) => D_DATA_IN(6), 
                           D_DATA_IN(5) => D_DATA_IN(5), D_DATA_IN(4) => 
                           D_DATA_IN(4), D_DATA_IN(3) => D_DATA_IN(3), 
                           D_DATA_IN(2) => D_DATA_IN(2), D_DATA_IN(1) => 
                           D_DATA_IN(1), D_DATA_IN(0) => D_DATA_IN(0), 
                           D_DATA_OUT(31) => D_DATA_OUT(31), D_DATA_OUT(30) => 
                           D_DATA_OUT(30), D_DATA_OUT(29) => D_DATA_OUT(29), 
                           D_DATA_OUT(28) => D_DATA_OUT(28), D_DATA_OUT(27) => 
                           D_DATA_OUT(27), D_DATA_OUT(26) => D_DATA_OUT(26), 
                           D_DATA_OUT(25) => D_DATA_OUT(25), D_DATA_OUT(24) => 
                           D_DATA_OUT(24), D_DATA_OUT(23) => D_DATA_OUT(23), 
                           D_DATA_OUT(22) => D_DATA_OUT(22), D_DATA_OUT(21) => 
                           D_DATA_OUT(21), D_DATA_OUT(20) => D_DATA_OUT(20), 
                           D_DATA_OUT(19) => D_DATA_OUT(19), D_DATA_OUT(18) => 
                           D_DATA_OUT(18), D_DATA_OUT(17) => D_DATA_OUT(17), 
                           D_DATA_OUT(16) => D_DATA_OUT(16), D_DATA_OUT(15) => 
                           D_DATA_OUT(15), D_DATA_OUT(14) => D_DATA_OUT(14), 
                           D_DATA_OUT(13) => D_DATA_OUT(13), D_DATA_OUT(12) => 
                           D_DATA_OUT(12), D_DATA_OUT(11) => D_DATA_OUT(11), 
                           D_DATA_OUT(10) => D_DATA_OUT(10), D_DATA_OUT(9) => 
                           D_DATA_OUT(9), D_DATA_OUT(8) => D_DATA_OUT(8), 
                           D_DATA_OUT(7) => D_DATA_OUT(7), D_DATA_OUT(6) => 
                           D_DATA_OUT(6), D_DATA_OUT(5) => D_DATA_OUT(5), 
                           D_DATA_OUT(4) => D_DATA_OUT(4), D_DATA_OUT(3) => 
                           D_DATA_OUT(3), D_DATA_OUT(2) => D_DATA_OUT(2), 
                           D_DATA_OUT(1) => D_DATA_OUT(1), D_DATA_OUT(0) => 
                           D_DATA_OUT(0), PC_IN(31) => I_ADDR_31_port, 
                           PC_IN(30) => I_ADDR_30_port, PC_IN(29) => 
                           I_ADDR_29_port, PC_IN(28) => I_ADDR_28_port, 
                           PC_IN(27) => I_ADDR_27_port, PC_IN(26) => 
                           I_ADDR_26_port, PC_IN(25) => I_ADDR_25_port, 
                           PC_IN(24) => I_ADDR_24_port, PC_IN(23) => 
                           I_ADDR_23_port, PC_IN(22) => I_ADDR_22_port, 
                           PC_IN(21) => I_ADDR_21_port, PC_IN(20) => 
                           I_ADDR_20_port, PC_IN(19) => I_ADDR_19_port, 
                           PC_IN(18) => I_ADDR_18_port, PC_IN(17) => 
                           I_ADDR_17_port, PC_IN(16) => I_ADDR_16_port, 
                           PC_IN(15) => I_ADDR_15_port, PC_IN(14) => 
                           I_ADDR_14_port, PC_IN(13) => I_ADDR_13_port, 
                           PC_IN(12) => I_ADDR_12_port, PC_IN(11) => 
                           I_ADDR_11_port, PC_IN(10) => I_ADDR_10_port, 
                           PC_IN(9) => I_ADDR_9_port, PC_IN(8) => I_ADDR_8_port
                           , PC_IN(7) => I_ADDR_7_port, PC_IN(6) => 
                           I_ADDR_6_port, PC_IN(5) => I_ADDR_5_port, PC_IN(4) 
                           => I_ADDR_4_port, PC_IN(3) => I_ADDR_3_port, 
                           PC_IN(2) => I_ADDR_2_port, PC_IN(1) => I_ADDR_1_port
                           , PC_IN(0) => I_ADDR_0_port, PC_BUS(31) => 
                           PC_BUS_31_port, PC_BUS(30) => PC_BUS_30_port, 
                           PC_BUS(29) => PC_BUS_29_port, PC_BUS(28) => 
                           PC_BUS_28_port, PC_BUS(27) => PC_BUS_27_port, 
                           PC_BUS(26) => PC_BUS_26_port, PC_BUS(25) => 
                           PC_BUS_25_port, PC_BUS(24) => PC_BUS_24_port, 
                           PC_BUS(23) => PC_BUS_23_port, PC_BUS(22) => 
                           PC_BUS_22_port, PC_BUS(21) => PC_BUS_21_port, 
                           PC_BUS(20) => PC_BUS_20_port, PC_BUS(19) => 
                           PC_BUS_19_port, PC_BUS(18) => PC_BUS_18_port, 
                           PC_BUS(17) => PC_BUS_17_port, PC_BUS(16) => 
                           PC_BUS_16_port, PC_BUS(15) => PC_BUS_15_port, 
                           PC_BUS(14) => PC_BUS_14_port, PC_BUS(13) => 
                           PC_BUS_13_port, PC_BUS(12) => PC_BUS_12_port, 
                           PC_BUS(11) => PC_BUS_11_port, PC_BUS(10) => 
                           PC_BUS_10_port, PC_BUS(9) => PC_BUS_9_port, 
                           PC_BUS(8) => PC_BUS_8_port, PC_BUS(7) => 
                           PC_BUS_7_port, PC_BUS(6) => PC_BUS_6_port, PC_BUS(5)
                           => PC_BUS_5_port, PC_BUS(4) => PC_BUS_4_port, 
                           PC_BUS(3) => PC_BUS_3_port, PC_BUS(2) => 
                           PC_BUS_2_port, PC_BUS(1) => PC_BUS_1_port, PC_BUS(0)
                           => PC_BUS_0_port);
   CU : dlx_cu port map( Clk => CLK, Rst => RST, IR_IN(31) => I_DATA(31), 
                           IR_IN(30) => I_DATA(30), IR_IN(29) => I_DATA(29), 
                           IR_IN(28) => I_DATA(28), IR_IN(27) => I_DATA(27), 
                           IR_IN(26) => I_DATA(26), IR_IN(25) => I_DATA(25), 
                           IR_IN(24) => I_DATA(24), IR_IN(23) => I_DATA(23), 
                           IR_IN(22) => I_DATA(22), IR_IN(21) => I_DATA(21), 
                           IR_IN(20) => I_DATA(20), IR_IN(19) => I_DATA(19), 
                           IR_IN(18) => I_DATA(18), IR_IN(17) => I_DATA(17), 
                           IR_IN(16) => I_DATA(16), IR_IN(15) => I_DATA(15), 
                           IR_IN(14) => I_DATA(14), IR_IN(13) => I_DATA(13), 
                           IR_IN(12) => I_DATA(12), IR_IN(11) => I_DATA(11), 
                           IR_IN(10) => I_DATA(10), IR_IN(9) => I_DATA(9), 
                           IR_IN(8) => I_DATA(8), IR_IN(7) => I_DATA(7), 
                           IR_IN(6) => I_DATA(6), IR_IN(5) => I_DATA(5), 
                           IR_IN(4) => I_DATA(4), IR_IN(3) => I_DATA(3), 
                           IR_IN(2) => I_DATA(2), IR_IN(1) => I_DATA(1), 
                           IR_IN(0) => I_DATA(0), IR_LATCH_EN => IR_LATCH_EN, 
                           NPC_LATCH_EN => NPC_LATCH_EN, RegA_LATCH_EN => 
                           RegA_LATCH_EN, RegB_LATCH_EN => RegB_LATCH_EN, 
                           RegIMM_LATCH_EN => RegIMM_LATCH_EN, SIGNED_IMM => 
                           SIGNED_IMM, MUXA_SEL => MUXA_SEL, MUXB_SEL => 
                           MUXB_SEL, ALU_OUTREG_EN => ALU_OUTREG_EN, EQ_COND =>
                           EQ_COND, IS_JUMP => IS_JUMP, ALU_OPCODE(0) => 
                           ALU_OPCODE_3_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_2_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_1_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_0_port, DRAM_WE => D_WR, LMD_LATCH_EN => 
                           D_RR, JUMP_EN => JUMP_EN, PC_LATCH_EN => PC_LATCH_EN
                           , IS_JAL => IS_JAL, WB_MUX_SEL => WB_MUX_SEL, RF_WE 
                           => RF_WE);

end SYN_DLX_RTL;
